// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
mH6KTQRQTa0hvT26hz7tvpeKtqMOdaNe4HtrFGk/RsNAIYrK4mV0OHpF/bnEJsKRKESCMYF3aNJb
uMJ5q5iDpFjS+5NqmImS+I10a7vyA4dRueglWrmPbkSRvhpEIkZgn+r5NAfBmibiQczqT48Q/NlJ
tSS2fFOpMRSm+DoWin1zbOwRiIoUXHgtRzBuYV01BO+pmSlGoptwSrK6D3uZL1gYBsP+4M7dALua
U/9YSk28rzCCJQXnFmvSysfMcnKur7cxjJFmButq+BIKWYeVwKVpfndO+3BKNm10CRvDWTbeD7m6
AeE/2ZcdQLK8nJt11HvEeS9IJoynQUgWo3WqUg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
xEq6AnyfUFnqivy55PsQPm5E26JO+X2D+jdPkRutgQD7WrlQmpUpLnGym+AOJ597qLKV9l4x6Z4H
G2jsPeXJh2E9iMzAI2Ry2wJWdWbqQZgqOzsjV6jgcxJe7H9aRdOO1Ct8mzmlsQ7BB2XrF+vTdcPz
uZ0VFDN2dSlko+X37nnPs4bdjs4530h+MyPA3SQgMAlweFsl/JU/5sudPq0aLVRUiL6wkTjGhMLX
jiHo/GM3BCq1DwMLbVEjXIE5+dnVO+gP2yZHFiDb3Yz3r7LVRfRfPycEc+MqLVhY+lp3r+2dVvsW
92aXgkSt6jEqs5UWvZEBnwp4+l8ztCALG8IRnjcWEQfWdInz4g6+hfgKdfOb0rnyp/c4GDosRaOb
BIEnq0gkf3am0uQ6FncSK9nNgyONnclMeftt5Hf9P+EHnIRGEdxFpmyeRUmPG88uSabcEtffJeVL
u0Qm+L1ysjTv5Wn73JR0k8Dm6zJclaMD+qnb7a+h71qy2HsDIGWxyXV9k/vGciR3unTOY+ATTPOH
9aZwI9/0UQm3f0bDDZYqJvBzmX++/S2co//mjRG4yG9j7QJVQYALGZtC+fGVoKwPIVFkoncDX8kw
vhd50DPKorMEotzSXhdVoOSJtlQ0EjPA+yLbv+AJX3gkH0d6YGBUOrrZtkrxg9b8yt1z6xYQRDgN
YddtPIBxEvwvhQ/dtzlYBeUXa7eX6/KzR9pTb9Ex35gBKVM/tCOSQds/CnU4mXX+Umcy/K9PVhKl
BrjeGWptarpzLrpxF6/i9KyQzZKrU7hcYXglFNBigLV9TcR13BX5D8QYTntcFPcXS99/4VtVKqkk
DPtkbYZdgTsWoY8dr3knh6uCBfywauFCmqs/ppMDLp63d3nB9juiTmXuh36bC1QCqGsnCmNSdqfx
cBzx/iqFosyf+kVd/bhkNS+9oXPZD6kglWiylOWL1MlCNUxyy7F6z09CPhZdZr0fLQziRvPntGc6
084ZZlYcZyc7oR2IZKDCKaeKQntSlOMthCsFUxDHJxr7QbECaHndG+Ulrr/vDrS32N31iBQHoo3u
YoP1Mjbyvvb/I+aTfqFEcST8wsZmkCN7iowqfk8h8ovzRyHR7YMpbMHavY5orbMAJq3QTLzHmTDF
9vw9/rc0XflRdF6jwkqwd6/UEoDrsr5hp6/z2GaxHR9Em1DdYSOybOelgWEnykaGDkUpVm2FbmLO
pppNC1q/XDt8v6jfQgY8iVoq3HyhxNjlWDic5MNlRVfkacAf7O1xT8pVw8K/WU+YKaU20qgM0QTR
0XGJixqnOZjJbxm+vDZYNW89B0TIVgxbgILSCElzYdTeUwrmAsp6RX6BX+2hZScI4FMSTS0OXlFr
W1Nfa8oZ6QDBhCQXcKbqJsSdQDgBTMIlTUlTILzzCH3sIs+76CFfT14oJB4/kqM71IWbcq+ajI49
NyT2xMpabsBMre7qE8aOq7qA1gLZyiYlJSnaCl3CuCJWUOCjQ8zKw7GpqKWnjoIsdXvVlZIyqkSk
qD7j81aYZduyf074k+/cZpNSv5uW+KRnlqAewQHztsmpYPg9QEkpglREZQ+F9jAeNaMD9W7ivxlE
yaHiIfo0QOoUQDlK8wTM5xAVE0tZSRr40dFLZndMBF5Yjlr90iTzSCRZOoveGe/89BmvnB5K0gtI
2td8BWwmkV0OoQz0XvQxUHpe2boZpCKsAxn8rpxVJxZGNqEjmJI5tNcVvSbozVjPsYMVaAfMh9h2
BNv4SlHOv0wKTVyL+ovFz+SXILBjUzEMev27xGQmBa6YvKGvafUlx3NM52W/Jp3jAw4zUSkwbnmc
80Z9Ofh1fq8iSpdAU0jxbDOn338/QgnEn7fkBJsGHwxvRUKOoQGKdYj8B2EPgEP8Sm7PCVAeNaBy
HNowIsm85AYyBnYTQ+W1jhpA46/GDFTLn1h/dZWC3eBEeJVaTFb6NZyfrSggLiB+0zqYk5M4cRf/
jHPGEUiNaA/Bee4yCLQp44bgRqCuAOwiJxCrtM7LEPqhux+KHzCnNYYHOwuvLSnbtFLHoK3EZaHx
vOD8rw2WjU3+SPqpcSeQdK+KPKxxSm8EAMsb08VlizR9C9vQ6AHcHPagckFXYzQMFHyvng1vvZjw
zBkE+e6I3Ik6WONNnZlF/hXxlUwmEq6UIQv3rH/D5t0MbBXO3oY1X046vJP5d2q7C8j7/JlekW+D
dbFuZEYseTwMi6Bx/0iH0Am9mOdvJxxs5RTxjjxN4TUGrIX9hZunIXPmtNTRy+47TcFZ2GVPKXK2
eMtuWzxGvMJoFtufun4Jcxd+wNzny75Wu5GC3k0NhJ6y7R5XOnDlfbH8u/IZMGp2KHIaGE7CZusE
OG3gVDvs80k4tyaem90FYBZDM5ZV5F/xURKIE7Qd+CRYfwhLTCUD17N5xgkuOgEni8LJjLJJ7e2E
iGbkZqICpE75ShduB1QX6pfMr6t2r69QNMomDadAkXy3N7DtNwBNbyLBrwbVWwYnw0pnduBAVaJ3
OwAVqzCVHC2M5gXOWI6t9ayQw3X/UTtSglgb1WhpyG6NIflno09Jgnjm6ylqnxb2ml/Jm6k/y4Fx
IvKUyNPRWhG7SWDXnO4aXKMl7IVSv3He9kGalWUljMtXrEw0yX/rw8vY39LJrgl+2TqXd7XyDTfG
E4w981zugxmrnxsSceoddB3CxGJdu/9ZSRYbQSfGCCO4PjJy0lLtd79ksIVoCrz/dOez1S9V4tEp
/08CK4ZcJoXvflaDb8gVKUCmhOnxi2jcJe4HweyZUezBOAFjMUwWQlYwZAWO+/Btqfmq0Q/0Vs/5
PUQUKpOyRe7lbuwcafNhWw/w42vCb2iopn523rdJb611Q5eG07fTWOUo9VXqbA9zggNjyj1TVbR0
x40A1Y/LyBSk/tCa79WquBV3zTATc+TNaeBifzcDb1l8wcUxL3a1HJ2BSgltW7H4NCZCD/Hgzgg4
iOTaxemWmilb7G/8e4bEnDF+9Gvt8i7GxgyA0eJWm0nGKXYaNAxUMR9v9s4ARPMqg9ZVgXlHahGS
K2+qWlxY1doNuRDj+ziJ+fXKan3gTbfbhqccUse79XkxTvc0kUXKzv5kZQJ9F82d/UI9tPtht2j8
xD5Aogn8lKVZnqTnPlkO8KGDxnZVC+YNOdj4/5VMDMMFynsq2FX6W5eApcGYYX/M9pQygcgqaD/j
qGZNKbnf0v+wen8s+YrGDGKBLAgDSfY58wKzpoLi1rJOs30b5laE2XCsjJO42uS1guZdBghJs3ey
G59g/H0ZAFEEiHkEJmKYbsJQxbkobDYiQzt9xNQoHup2WrlJCL1hMtgPiMYODXkxjeUMEbC+P5jb
J2QSQS77kcOgH1XsWf74/9Hhcd4eikDElY+VRbKXL/Tgr99Jm17Zip2Upm26fReKRKvt9W0VfAKB
zzD4sCNl7O6gf/O1YtA7qhE/NJnEKm+qyo8m6fm8i+Z5g63Rnih28d6Tye3xpJaGoEFzJ0ebYhVn
uW4MOzqUMy3jRSKYQLaoI7X/Rv019TsB1ShuPoEH/OTso6jVxtyOYP+v8tRrmL9N94I2yB7HQ5nw
jq1lXJBQcDH0mJnhBp9Ty4B2iGdVLox90SGipv2cPimhLkFu7spnFP26hqi7xTeVnJdUVgZRpTcS
ozAZMJ03nl2jXNrzR7OQ7CSyckPMGZ94nf2fFcdlJ3Ntvm2LQPpRg6JP9JSDzfoezVNGOmp5q8gE
u+QJotmzB6njRxxiwxenhay7rufm65rL1hVkXhv0WVkFUzX27OncBmgHmU2c1J+W3XfBCxa8iUE5
jqOzgDSimb3q5JbEYNbFuzqacWn1W6kQ2L5EaWycD6qBsulixwdWn4fbKbU8xDzddOewXzfUSDNW
WZmbfLduWGIGDoFPiVZAhcRlo+F4Xgw1JFzPbmpoWtUMjCLQy2ZYUaKbccOzLkg7MxxA384V/7FW
UvlnFHpJ97jDg4pmrYS3zKhCR1YW/7S/bTd6Mf1ERmriYwiwHuef3wuK7CzaqctpdeL4kcXv0bAz
wowIPsyEVJJfuQpscaXIga/NbV0PBfqClzVi0tHBi/D5clkm7mZ7oNYaZ7bWzphmePqL3mL3br5e
CAlqy1Igl90QQXXBb7obPybxTjgIGEdqngIOlV9EDEEJeK7Kc4mJNu0rW0DI4RvEqraGkqoJHfNl
Phc7DEB+j9te2qExX7W0MCI1w0mjvlGKp7LC+7JKx9oGJ1TSXVkocjKAXXMo7u4NTKN+EQyjGFq0
V6i5zcg/PAxkSHMGruFx0Q7PIt+2aRfOy9xuHKQXf8t/aFYnhqk1vljSQYT5QWLxCtnIvfabt7n5
MQUvi3K6jks6hg8BufllQMttT+ueQQKIlNw6jYqb2kYmVt2UUp+6Y2kTqVSc6+2pJjVkV+NfWBiC
8qN0GXfkWS3BJA4TbuuLq97AP5PhL+ot8QxK42uMzN7jjGYnMCnSWNPVnTM0WG2qElKoec298kgN
Q8JzJ4q9XgoKNAf0pyWdlv5T7oNLfNRARP21hZJHl/LHBISG0TBpIwDLV4yyPAq3g0d/oId6COPu
HTQrHMjApkCpHgmeDV1jkiv1NFkoOeLzeJNjIqRvYw3nIatpn2Z1CIybvWfXoLSgl1fO30MvhF7s
AXlIONXHDuIs/xkIMVbPSVvZieNn66GqOk8dkpMfmiPZENo/1U/RdV75vwYURRR7h1eyLgbnXz+w
C3ygSS8AXYZIvMjXmDEx0W6fAoaxFd2nvu7R7VNEE5sWmPoGPGcud0vBQCDRp643FDm1jF0qh93s
35QdqIQESKYmKu/9wYX5bublIy36BnrKJdSiUUJwbI9jmkU3wAOlWoD151HzXFP36LM9JoCMTata
VYJk0PWGUE91D6Pkep5FX2NG6IM4KBDm+kHGZfsnegicEDP64XQD9sp191/g5dYFAp3wNsR4v8tt
6KoVWq6qnU24QxUHcRzUtdTqgZbdX14xX97Y74NVVy5YMLXPovm0fCPWeI5kHN0fTKnAfRVqZ046
Tn8rIm/b63OPPOqM9HjctrLIi0JKjlJn2+WQtL9MMSTqk/0PcuwiIKzKSDFfuQ1BQEyWwB/A9cjO
vZlAPI8LkzazHjYny2OYMkjLmhiPqT67wViKgwlK05nSlj8MJYwjpFADl6ZVCTXym1YU81IF0zYF
7c+pCs9aX8WIXUuV2cFxf0tWv5gB4SymjnpqhbZwADLVNTO08sOT1U6ZJgwsoXX5Prx4Hv3ZtZay
J0PLC5i1T9cTpuJRqczotsQS0u5PmMRJw2ZbplIgv4y3/weUi0fAx30XLQXgb+lbnVf0M3DF/cjx
WMqY9S7nOMRB0gFtK9Um6XXADRFEDPs5aB90+yZDv9DRWYKhYMUYyabf1wHYhGJzt+Yey7gakjGl
0Tud4Qa4nnCP8xWHNHiN61Ye086oIBZodmGUMS1EfMQZkybTSkWQsDCO/aNXAo/aNJsnAoZW2Zuf
ZFcFmlYAc17tBS8KXaJaUibb3kfcDrQYeP85Hejsa8ULHZBHoKPrbQiRoEiCdFgTE4ELr7NSS2su
QbnVQUpIR/Z8POBbnXpVYMKQdXq7Xj4H0WT0sS5W0xEKCVH3gpXtUdfhtfJStLc74P97nARMtVUv
QCBpkY0BYrxfMnjpvMwJIjZr0BZqbQdfNIpLSEJup3nUDbDEu80aT8I7nTvopMp8ch9ymq3E8bMy
9DcEgcpdGLHDCGG2wV0mnwN0y4hQIRfdm1pEVE5ynQp1AAveNYKzDtysXgeK8QFcn5qGVCRk79+x
huRoZShwJAGLC4GLHUcTwSdW0dYchlm9ft23Z7sCK6NdgvbDjyZxr4P8g406Rayh3Dv95v36GRTO
t2TbicoV1iVT9OR4gCgME+lB6saaD1HUxzkDxU9abzpCkIyFzjTFkPco0kEo/tV2Gm3MJTOU7p9e
FoASbQkUKqWQhhDx8e5JMB3MRdid7rA17blU+UXW1mqW0EiH89S67m6eWd3NyhRuSP+KS8Almybi
f3BYI25t9mtL1KQd9TnmRWjJFBJabSyyH8MRMDtclp/zEJ4EOEQw7Ddayil+VJgg2SdCLkfRYzN4
erRI4qD9A6+xOtZ9xjGBvZ125aLH1ixV9BGW8eJpqzkep7TMsKv2EApQG0aounPWIPsbriqs1ZKt
mGt36dq+c7DwWBIn+uSW64rtosf8GMDt8PuOqESjpVhc7d56kguYKhvPJ65JxFPPH6QLnQCrjKVk
4gPpoGtVA48cuvkuD96rby+HfJ8V1jQj+41AHGCmcotq5t9DfBvyGtlSVIgslnD2isSwVJSyGvXC
kV+KELFgqu1YoJoLrfPFzxb0cQ/ztS7n1Z3G0mVfWm4uNB5qf2opIC7l7YWb8/ChTguYfrkHuKc0
nFaWpWxwPbm/Bfy9IVWri7huX7Kb22v9Zihh3w8eTicirgv9xkiSNubPuHH9mmLj8h5QR/HG3yq9
F2IKzghhq5mr89neBRiL+m2KzSbmpHbZpWPsgG+ffASE/r4GT4tFPnByqywqn8bO+KjFKGlp6pOt
kMHTjGrJZAh/kOd2zw0oukErbe5qLeihpgz71elcwUgXTc3eRulk1HEW3KFYudvf94+m/N808qWd
PusvwpJrRUD4Wniqb4/oOG3tWsf3am4MFgAm5LH9/zpwo86uFJ5y3W6ycTug5R/4xD3auStBnJpK
QeLEVhb/zBB7ZA4QABPAkazRRz3Y4EJFmv7worP5L3L4SbHZVPncp1dK8owNeZzfmbVugB5hBAlX
+ijzmj3XoyEBWzkX7JZYNhEl5eouYcFsFpQJiUlkNRnsaurQeBqg9OzfhRrdU92C0iJmajvWL25h
w7Ew/aqacw2m0nGS2KExL99fUPRCLyx6neVmIQiKW9zUbf8yBaCPsCSg+9NTVkBmQXz8LcDhHayv
90jhTb/l+K315C9sdnVm8v6k33AIiUQ2hGEJDUG1rTwEMjW6e1R3Sd8L1VJZzXp7/hG/xuVhrIYh
JuOfOyjkkjnEuWSmFu+RIjVPzgtjUJVCvcmzIc/OLMIqoS7IXvWxjeZDQ8+XM4fOcx66g6v31LHF
KUbAnyfsuLfMScalW1iRvhyZxs226g9D3BRLEuTwBp4mVn/lhxt8kLG/OM2T+LC4L4MC0fqqkSu/
oy7q/s5Yivwr9dvPzbrzItTPas2yQSB7ioushTfw5I1yS8z2CDlQjLELTB9S99YpMwxDyuR0wI9/
VT03a1iJPMkH+pUCnBHYHv+1bXzFVds5BP15kdjPS4BKI4ahqxS6/CWMjdECYsW4/MwjMQjgckGR
CsO6U9ZzSwWs42vYhWFVQQ1+/PSgWMlgHhz3EvCui3oM3r+cKBZA2UJZizjl6QHRUocwqFnLWsnr
xnoaZ4UPFWrNs/XXvLuObRDZMq+vrobRZmj0pk+BQazFQoKYbCjYHVaYV5xEXMuTJlay4hEfhprG
SEZS3clBQ8XMJr2QufOa+VDtgo8O84YPKusqRpzeVZznEGdfu0UTy9ank1wbh4rr3A8lL2umra8Y
MYefnVOV74Dfl74ooFXEkZbDRUpM+0iKp9ab7X3QbxamV761KGv9LY3h+Au4XzrIA7yeztna9mPe
JRc+z1g/zTnSIcXF5SLhLpT6ZHyZF1MjXvhqtKPOkPJWaKPbP6dS6KSeoBr93Iq/JMgiehk1w3L2
3a++HhwUDEUyKFIRXq5CuE6gf5thfQql6nWrWRUeUM/HdVfwlqt9gT4nBd9VtD59bKeJ9/vh1ZHM
tZB4z019pbG+M/znHv1YGQx19drzjmJ6TQdxwWKfRhHbsZ5B51L/zB9ouE2b0ATYOE5sboGvCdaa
PzjkWx/Ho6abXL0MGHBHiocu1Dmkc/q/VK2Yii2Gya9iqBVmtXtCyzlPH+2NCUT1eDv7Pc1bvNse
KyAeYcLLojjn2+jtNw1BNWJ6/ZV9s9x30yOfwpvliEZD4Q9TL0L5Pc+9OUPtNxgh+rY4YzdY1O6R
Wt29WuiXzGWPZUnzrTVXtNWNDuIWrZ4R2/IeC2I0hvVTyBb+0hC5pKrKyvfv+R+wQafkRA74kDUk
CHAMo7JdtrelWPCVytQcyftOGu4+SuPzgtG3quswf9gIAo3fxSvrXpsDESXEOHc28OCq5mlwqAl+
4Ng8lvEzW7vmcGgVmORh8TEUeEC/uV7HFE2v347HZ5V2HpfLpmK2UrlpNqKQIUrlBG6o0747hlfB
nNKzTAYMP0XPzhT2WXHzzAOY8VhzA9YqIlQBL6HiBziXaNJzOIjhAj8EBxepCSk20l7jqK/ELkKM
x0Un5OYjdAEYhWPGRaiS5feSfyCIlyYObe1WVmNv8jXKnX2vv7hZdFxvrplFFQVVgybAqq2LDSxc
JAizyOyHoANfcVoZkUVVMIIBCpWV9aHf9HQ2rwQsuwcs3M6gryhS5YmW2GGdxEWim+xIVFdTvsXF
LCj18jQ3VsXFur4Jv5QG9DBW7+hNdTQih1phhqIyptGL9jHO9aX+EevSaRNGmYzkIOumN+/HBm60
Td16EfKwTnqLCbsJY30txCkdb1ZEYAqbdbqiNaPkpAhyYC2GG9GWiizyN2zkPsgs4r7N+Eaiqkrm
74mKt8D7R64uojfHUMHC/Ha08lL0eAkRdmRn2sOd91CoCD3aDeq9X74JP5RIUqctAa/j2uTztAzG
MRUC+ALadb3Dl1wI2LetZhjH2qCMIkHsNufSt5pgq7p8MactQ6JuIPDEV15V8s3FMhumL6hFiiYs
zKrOhVm/sue/Jv4sNoxaqjrEsIkZ91ELoIEVc1Jf6B/N/KBAz24FU+vR7I3OQCAlkbiyHI4C67Dm
dI0MPLeK9JqZ8ocPTwujv7f8KzoqY9nY/NKuDcRSm77BQzRNwG1CLndPsafPG4JcGetgnF/PJZLg
t788unGzZ9I6NOzh5xqRs497MJk1a9CzgvMgAU2UCoj6cU0zVbqGKLcYwsNhCsL+wLYrjsXirz4k
Yb2yBXSF6FLEt40BUq4Xvr21K+lVcbb7ruUGtj9weudnTDCoDx9C7F2hz2crYmy4vXVOys8OGdRU
OS/vS/NR4IgvQCwfdqSoA2EpadukcDhV6BpDdZlam6biXFpKDH7ZlAEE/kSIqUiDylyRO7yar9kZ
xMZOhSnipohWEj93vZFeaXqomGcmCf9M+bbov8YfsuQ0MuR/iLB6x8IF6JZV8i3axsgDIreLD+ox
BuvQrDOn6ClxRsgXRTVh1AGItUESKvQIWxcFSwkP935qYN8S+8QCzFUCrW7nIuISnCmPognismzL
8TZ92+U0PhaZtzOyDX5F60DWzNaJ2EbbJL81WH2VK86iqiXNftGnbpLVYrZYGDe0u0mfH8VtbtDr
v18f0TesTCc3uwQfOt+rcquzbAqUtqIRQ3eAKns4sFsOvdO9oO0YI8PCFC/cFLQ4Upc6uwpF2rvS
IKh+lBTK0h9m7PxTVN9f3BSeeKS4BAfV2CIedtwYJjygarAV1Gand6PPKIt+SxNWguHp0XwhKm/D
W+HVCE0oK82R6exOeKAZY84gzfSJFJG8v8+UT/x2dAemk6Efcx10iof1pSMqFG9eG4EhWql02+QB
8SPJ4wYCzKrgg1SpUqU2eiuJFUbUmhGUL0Kkglcru7FwJ3IZBO0scpGtVJ1lULz3zXGzwEda1Cc3
3LcxxxNDuvJdiw18P5jEU0ckBT+KS1Ek0kagAF91GieSFPrhcUC/ShgolUz+p8fa0bmBLwNA+ORN
b0iCB3foxYaG/UJdTP8s+cu2ma/qDAGc3sSVgxm0+Lqo2cA8curnKYJpfdPaHJxot1Tp87Dpsgjc
wG6k8Z47rxQSK/DHg3ALyE7VTKmV4UMZ2Fa5XimdoBn9fTqjWFzz4RqikRm+Qx7hpzTM/lWkgyoT
OXP9EwbVJeLrlheYbOPsGOIGY3tDW+eY4TvMPTKF0bL3/jLoH8xurfs8w0EN4VIPE17GItRiWN+x
P9uAC4GuBEYn2kGCm1Kl2WACiJmBTnwN0VYm1kuS3NHPbGiyT272DiZsZVQrI1AYGxFdaBBg148Q
CIFtgWNvujiODLzdBpGDdX9kYzQAFsGl940x7efxxzIsZXEtfkc1Y+EEq6pIEFBHgUqAa/IXxhLd
jaUMWmyPIpqZ98cwi+y5+vX6ou9Vo8CE1mbAV5A+KgR/VrEG20cIwt6Url1cNYNUjT4LHbcyx650
f0TT651OChj4YUC693AuXp/IJi3GhNsLF59kyImBHoYrUHLuqdSQUxtrC7exEt6N+8/mRwhhCYsK
PnLOnU1exJiL68c1JmNuZndvkaw5C6OFF7X48c2lAc+qHAsokpH/7/61ZDpGNR2sNY67MVplkf0j
qBy3s1yGGG6DWIhIQm6qdYxIsyiFFYuvFZn+WtVzdGfRDSZYHWfYsmbXkiix1+2ZzLEY0UFatT0Z
fOPU1ChcQWtPksZyMr5IjfnDP2QhOaHCBnmzxFE2JL7rpZGCE+w2QVNFUEuyGfVf/68a5MNZUMUh
MGOiJsd1d21MY70ovCTQnoI1lj8J9wzTrLP1F8JtK/iwXwPifFGhX/s6zKw688hrF6YnlBPE5J3o
MpMoWMYpWr5Emny3fL6ELp2JyyFOU7ntBbqAJXwZJzkvDBMBtMgvOcO4eDB6MZ/3nv2jOp3hB5mm
5Dqt8Zhq34TzYx9mXlFAZyqS4AObuNCZwgjgYyTmXtw4nlHzFUDieCuQM8w+uWpnTDMhndSwrRjE
2DCS1uxZF981p2Zhn3bt69rlMfskbSdRfP1zICkK6NncgG34OkS7OsQ3VMSRmAO250BeAub5005I
XBZa2hG4aT8uBDVA0S6VluTiVil1Bvlxbm8tTohRXMKzxEmvEm7IPScQP2WWzA8aWqgqqtWpx/Hy
CeoRyaq9gtKkB3Vnk07q6BafRWPFo/AwmJUPuxf9+jC8TAJLwkg78qRzUbIOFUYm4sCHrHU7W8yp
DL101r9yTqHnHcRQseNowOO2nH/ZWCs/vRUg8uGr7XJTuei9JTIpdFi3/G8cAEnwfxn/ptZkfHrF
C8tR8W4bgveKFOHDtH9KOWZq+rmIjPoPO4Aq+KxXtoZ7EXO0upOBmwTStBzqV98YwFAOGrCloWQj
yFj4zaJXeDJk3pueDXkD0+h8Cy+X8e619w3VrZGUXT9vLnTrKdJdkGVKp6ih1s31PgBFVOArKyYI
Ci0caXVX63Z+iF1IAKnqoVxGCJOeQpIQpPcDQMuwuK+hHNZnz2KTQ+hSB35wBq3C/H3eRuCFfiLv
fGnmCt48ZYHigLxvsyQ/yRlzjnhX8STzPg+Evo3UvIYL4rwz+U+gYLxbtXbckfTUA9EYN4lzj/Ri
zKeczSOUgmesM2PfwASH2z1+zLQv5K6ThpXIjH9uKM2q+LtsJ2mtof4xdnCFi8wS6z5AFmYvzt7n
gPdVkOOfBeehuM7mkb3xwCUeQf1tgEzR1NXFVacxedc88mQQN6HnfEQOjBRHHVirHBfWM85SlhGY
Op0SEmbwJXskJNB0kA6sejN/xX7EST0sphErOQRab6DJqymQakDssri77z+TK+BLeAW+xgfqHMpT
9XkXi8nEeHWqf9rEcRHNbyGlDDTPzwIoNeLyUzVce90/6zN+jf5vbp+/Ea1uuRXZtR/ukGC0wMHq
iD4+TOcCivqQNxLuuubgt1UFkD6x2ocN3/jalYTvMyBuahKTRJO7a7Ui1FDhzsGdtVsWs1q0qnU+
QW54ZWvI6WRSFlY6MpLxICreC1xyDq09QQEHiIuc0xJ8c+MP+bN/FRGFyqL19Db7fF5HggqmbJiE
RMe5uzgJQy4bpz8NAVlEORkv7ZctU2sYjt+JWHaui7hhUqhjQ/jsyzVDLBJAYC8hTkkh4NRuUFMP
fpPivkClOWO+z2E20H6CXFij0VvD4RsAzU8cnwqD79ZIVN59QR8x++NGgoQsfG8GUuNQLDavbN79
5AtVCGKeWQF/pF+OESOBOc9akamxU6OOQA7D6h2FkwoyuMYAvZxWp32qaHZlMdMt1b+WSg8oWwkv
H6a+ZMoIMHofkEwJ+r8sr/dOdyUGIDoQ2lRz3FvGFqrgxar9KG2Pc/xMpjwszDJ4wUtYYC/Ho6za
kNKg/4znU7Kw71FgnwU0+y5RFA0TCiKMaGX+0g6oD8Nj+Cjm6IvSoNTnbd0yZO1EQQdLB+PLfwW+
myz8DofDJAr0yBJ74s+y3rJvqy3am5tSFa6QFxgR0ARKfx8fx6M6/OZwHmNTjqbuO5K8D/imfppt
UWJjJShFhWGnoKRWfbMki/thC136c2gsiABq48KQS5kzBDtCYnSfvJohdwa9D1RF0JUztFIluRE+
N0nKq/MzIUf+ND5bamS8Ji/z4OBPyajMreC253BbowM/WR9l2f0grsdBXbw21KmAS7Y7T4RhWLQu
DafRUbpaHihJfF2tRt5TVlFL0wAe12gOv0BqOSNugeGJQ2VfgVy26SOrhQ/477ph2TcOdj6D81Bi
E4CHcH49J20d2wGiFvXOGoki3Csu1TPTSC2IMbrf/Q25Lq1QRIRUJzsuTHW8KoiMuD+L45yTcD2k
vz1Zd38IzJe4zyp02THrkxsI7UZL3z9KmTU204HVqEkaKxu8YPbPN5hgJOcv+wu9bja6ir7v3C1B
LK+32r1JBGo2ymav09i+DcshUgYKD41cLmRPH3Mxp6l+NA/snMEuZYSy4+wsUWfyT/KodyDGY7Cl
RN28c5tmJx/TB++0+M6kiMku3DChBmwTqyyrMP7fc5eaQCJLmI4+x+kaPnfeJAW894PVt60DlceA
RIuvsCsdzqxLAi+OROKV+iKOD+Zjv6VlLzcTdu+K9IAobkKQor4e58gp+cZX4re78qOxVpT27gyX
HtLYYn4gbtSFlLAZSoMzPJSHAPI/e0VK2JqC0Mz8if8xYjVGBgGxTQJwz/NEQqWwilu6TxRMn/S8
Kk5TIKnJZuBZMH7D8yGF6atwkAGS0g0uKw+fW+CBkcRZ7qUO7T/V2Zu7Hnkhxl4LLuCdkZEsuS3S
pg9EphUhFYbyL6WAUoe36gyebrQJVn24W+Ee9IR/kSKIGtrP0LoT/JAINkmw6+gQGXv7lW3l0ruj
v3APN0z9Uulm29+gfgm2Tjg799n6yqCO1nIspZI3bnMwaBgmCGSLYRdUVIrdBP8OMFUDi3Tp4S04
xvgJ/4LMzz35u9G58/2Z1cGQmaU4N1s0bhWfiv6XA764l9WpNnWoRf9N7xZOqBU/P/tPWHjCvrpx
O6gmySWu4YXv3lBq/ZMvLuvXCbF03fx4BkbkL5hSidG/fOOpfRLWOfHHLCd38Tx7cHGry6dQmK8b
rC3FFtuUj454H04oxFjS2s57FHf9bPYLWzaDJpGQL5BTJxz/0HgrwfIKck+3FMj2Zzp68jXU7n3x
Zetu6bx5sr7F+3gpHqOwPQdkYN/6QhvWp6Z6PyrnTb39ROPYfk4a+nPDqeqKWu/9yILA6mieR+G3
qzsHn9kNeL1nXCuPx4g/NxevBwDdt0yRTd7eV0GLyxlzAZIGq4mj7DjUOVKzrPUgg7lj1rZWIhlk
0411/n7GW/Z7udQrhbau3y8l8TiIZFn4WFj9QoywyAvibNNZ9q0YCBCSt1udeYfR7SoaO4hOuJE4
cxFlf3AmnwwKzmcn0Qz3kXQoSR3p+0wHHlSJPFCewssGwnji8ew0IF7aLgO1jrKesinQrgLX0VB0
pTjs69WLCXffG2bjr9D7+1wJcBHfy+OvjmCTuy2i7rHNBJLXw+Zz6zVKypYXSsQUkn5qcezzrWzD
WzVSpLFHXMJDiEy35Q5nn4BFEDwaf9N3T4eRHCwacdvI6xkPR0Il1Hnof9A9uvmHvmOf7V9A7vn8
gqBWo9EvmywnDR8B+t5/q/SL8kAYmuIIIn1AjOq5vzTE7MKE8FPzDgcG/QwneAmDXQ6fq6e3OliZ
3rxf5Bcn2zcNP8ODhF2M4lNWksodj7f7NCPdq0usQEDPBG/j8KwqGfYqeejqXLjYaQT/PdUZ+rWt
JQvJcmvq0AL7mZSumvhg6NAOCYzmtt2cKapzpIkxE/CGS+KnNXhAte/9uhtdeCIeA4N24gyb7est
vFpV+2KrOxvg1adgdfuV+zZRJXk2AsA/FupeZVtqYtOwUdHc4JLxb53G/AzLmuu8IADx3M5Fm222
1HE+wPeXTf0OnRHyS/cl1Xq970UMS11PLy4MqaU27gouZbRd9ozGonKBvOqu/Dmb6kE/6pRcVmqG
tScymljuQhWfJeCUOYsJg/BO90B7tpZg/jkQsWch5erqG/4GqaDMiW2ua4qPBu+MEkr9agZiWN2A
nfyRYbZOW1rQk1qSTn3GuQffYDAGLs5EImXZOOA5TiKDi1oh1u7efflrIX9+xS0wmb+BVmY+H2WP
+XH5AyVuZb6zrKQdOKqvddA1XGyUN72BOC+9aCqcO3rnG6qtLk9Eh5r42FXUDK6PJxvVcWAwJTqe
D41eiM6V0qOmNrU3uQG5CzvehXQ87QdAsj3QMYf+QMp55tAdiVdyLNUcnXmoH4zSaBV/uutEz5k3
m1fD/ZAe7st3JWJMZSbTKQsGqNWU6ctz9hYjLRu57HGwZM2+5VOlEvaWkYW7ej1JMzn+EUecx20G
07lBKqGp0l6Ca/31Yga+wcRERC5T1qaRU5CotDI56d7XngXmLy2x7HbdcLsug3rgnqm4CwLIk1up
PE3VTZ/Y3pqYULGSuRNd6S0Fyrgd0esEO52Vyt36AOlG/vU80fVsIdCK+rIC2Y1c4kPMRmYUneYG
3P/vRn/N5gVLpAxSYZeolww/pzJ9fgpiL57VTHtZRV/dORu7W+2N57S0Fhvi3nsmeVs+9gQfCe9U
30jkokt7HqNisXE14t8IM8yev8ZPAriKxmArPtD6m87im8k4f6WsRqBzj5mAaiPvmdEp+B9jguUY
NG4ENUiLlAiUMnZ8U2hqPn9HSxwWa6bAiMx9AjC9bF67zj+cVIXkHFEAZLs5M8URok8cS0rc2gPs
eBum/nyWcSwgUnQFwdVkFlSBX0XBh78oNVx4y/hefKb6VWYWvKbDiFN+l0I0V4mR6574TOFVQInK
jdF1HUyofjBQnXZRYJCaKFWtm+RE3B51jbXlkGokihWTgfhzFdeZUZr7VQXx2T1jvEjBIVVUxELN
Plf5cTAMjQDwQxXSJ2FNsATUjX06BMDhGwkQNZaAI4hsvMXKwhR8kUf0kW5/bDNoLrpN6E++0BFd
mKFa6F/VMh4R5MGhtvlLq6w8e+8JnfihhxTLNTGXX4XmEuOktz83juVI6ZW4xtgwLm23/Fj5R38C
cRliY/rEng+1BPajdS5eS4EoOscuH5c1lE8qHoMIm1iU9f1T2dHvvAO3WtA09fz6o7p2FMwDIvFz
vC8aZVJRYkjNXdvRGZ5BwJpo/5iZSEVAibyKDACLEqfVIfcRdOGO7964KadRYkS+9mhu4ScfEwzl
SQIxIBcwn5snsuki4NwRMb/kS0nJ3XI986akKJegaWY2+OtQGawQUrRBH7SG7FStsvL1e2cTbLjK
z3DhxUtHgWE+lS5x6H9SG2nfAbKKrqjn0hLGKhgekuVoRI4V3Qrq3BDsQRk+liCDI/o0+YLsDYzb
69eT5W+Miwe9TwmoCE+BYYC25t2WSs30MQlTQwNfAOSnrHKtWEWw/IG1gmboR5eXu2rEBEU+LvzC
kCzU+jroSKZV7+BB2joBCJVxuU2HgbuM75MTuUDQ7I4XZWFqiHCXBu1oexb4bcpeACHPDOUJvBBb
OaVKLMu9JWO5zar68zay1AlA2ZOc8/FlgvLNARXcohnr85CjNahiI5Z0fgjllkFybHDOpbesvwyX
jV1hqneAuyIKliG1Cg+0bohaNmWXTNhFxWLSmjkGtgRkrUuC2A1lDl1dUcXkG1Y3hIqlHs9EKUdz
oEeYUrvtjo7Py17O27Ddv1cr/8iffIS7/87FDBEiidM4c5USuZCQIhW3TgCI/1WGSZufVXZahzfN
fFntEUJlHiXew/H42Rno4pgmw55CVl1+T7O6LUB2UtfSd0eOHI3Szjqgj0IyosSn4QZsKLx75BdY
FDNxhmys838wYrLHwrtdufKY/dQjk6GR5tEGcWo8FLKjCPFbf6m1CzkT2LrSggFXneo43pU+wo7r
Ex/iIBpaCciNtzKlnWMG04f65OOWon9RnKu7pP6st98DB6mcZHy87ieblTQ0hzUbKQknXtw04Pnp
2GXSes4GFQgUdO1zzQpy+5ytzjSYfTC5rHUtq+RXomHhW9yT6uMOwfBrki2OoFtyiTrNalQyA6PQ
3F0p6fs7BjEAinUI8SPd0L24X9Uy4vy5uNQy89TQyYgpsq1gSdmShTxEFN6MwTodhey+2J/6PGwg
A21l4AlxRjeN14RBNQ4leECt+22SFVzuCcIFuSg2aP7V+ctYk85ZMeOk/Og+mPnXc5J5rNQYBBW9
ixTGdLNmS2OSrgoANnt3EiYUne9AfePpNdx3rKkZx/vJIECeUnCY14sjdKC7Af8QXMzTFjAQdI4A
dsw8PUu/h0hWfinUEtUiDqc5FzxysJVr0+DjWQtvWK3FFWV37aJEJjdxPHFfzFqY7xC1+T6jaCB2
DrJvtzrx332spZd/wFpiqGyeq/kszgMEG3EFl7AB0YlmDlHHsaMXHbuTEAKuMQL+E+ooOSImteKQ
pQbS4F8ccX5V00EuEekC0sG1nFB0WCq+CsMxryiMcpRRT5lOZd8ZHbzGm2QVC0/D/wVgrx5DYlwd
jmQV7GRPerjqcK6LN2L90aWEpJDPYwLRQzvoQnEdqAEzpksTc5XRKMqzzUhCRwli6wtAxiT690bB
hrIYz+mEdwbEXOSelknvAh+EoNOfwGgMyMsg90DaPNqs8QqNYI/YcN4+Gz6K0dVKNpEijcwYKjho
4f5WD35MCGrez09ktSgeeEULKwnzpZHipHPA2dgOvRKFEYuZF44GX+91J2y8TNwntGFWCuXfLgKL
3A+sPmBL2F5KyBtG6BA/a1OsTZUA7Y2ovlAMTYo+S02Zcluz0CKwX58RbtfvdU0oiwPLIMSE+gtW
7FZLEI9QgUVxMkZzuKdDSenLnHTtU/Tou6dMuqTpHHdyUL1tcwrkqKmz+0t1q+BN1TjQP6Z8BTnL
dOXeN8Tv5RRVHzU4UqQkQOmlKxfy5IYTUTJE17cKdnd+11ZrekCfecJUeUPucijuI8wZj+lVaszz
Z6kZO74qhGSBcnJ6KhOCzPJEQLJZ1V0QRx/upco6QKThvJ7FCdg4qbgJldraFnZAAP0diHWvqJag
Eip62Yg34yKE2/Ui+rW82USNBZv9UzHVuciV6OhzLnsbeSO3BajTLS8/OQcCzAkQdQAOmPj8q3BV
Lny4zQR7x6FaYAhggm+MTDYxbMUg0Q3kGJUI0TTfBwZUxmJT25E3EroGti/U5w1K8vIAHvGFHeON
Zf3QL/4b24RddUUUghksyCPERgTI4IHHu8kX0oQYLUWR8clkVVit+zsHVCfGVzghI6OKRLdVMWB9
Shz/nWWiKzkOSWr7wqUHwk14vicxrR3nCcgZnlecyl5NjRkqmzULQHqSD7/DDDoXywCLAER91KN3
G1kC3u19bhV6UD+TGnRXB6iWSYjfRqwRZ4jzQ0iKcrnBjbefb1OGLpVQ659WCi4ih8E7OSaaq0wb
js8aqoAJ9yRZsg5qArHhd83SHUaf6Jp/JEkhbXyl2r2fvIndpLa4sdSbMMwGACAHWq9XjLTWQ3W/
C2KjwJWAeACUGrrYUrEqoRxSkiRNm+ZE/y3ddNh5oqm9ygOs069ifpTfp2eAF5+1n/9V52LVvTnW
+wxJUDxok+ik5ErPCpQOLdl+yNOValF81BzVyWnLevJ5wDgIEpSWtoeKCDMZx94fpBRqQqwirpFw
eMC2RPoK8DmNUaU+72BwWZfyf2Ropr6Bm0S7yGeqRlIV6PNW5D8IzRJ4v0BDQ80lMQy7cBqS2mnZ
i8/sjAtuzVSQ1pRiGbxiArxSE//J9zJ4kvJPMBN0nHSFHxTz1ZpOUcBE0gNmKxayBw3J2pL7iNQW
6xSITJI8qHx4CJVzLi5csy0PLamdjkAY+RU/TmzBamplU5LYSZrSSq8ubP2/xFAe+oxcDrxUynUw
XVMmBrKKVyDltUvXghE48JGzJ0S3Rsxu9iLfBnUZ2Zmcpa5ASfInbiqJMKMRXZVLaHBNhgfs/RKi
6UD3MVajqKaA0ltoFdugIkS7a8nxGNSLJKeOmbxDBhIWPDs6bP99Nz3UI1YxORFroHauJ1nX+AgM
nCL3qhggIVch+3uz4riQFHRIGWn93gd3XJPV1IBTZYobkr4hI9KVB0spzoOaeKoxxx87v3Lp1Caa
SO08WePEvtb0CVdm+f+tSvggiQ1HIVpWiz45DygzhPeFEjMSh7Psj+RdOcJO7PbV2zYWrj1oXqiA
APYVIWqCaDae8G0sVJOnNa8ROHMLQJRAKj5krdQE1KGLSSQqriOr+0ECrndjGlE91A+WQD/8hgAs
qm+IAkdNjsQmpCKHU8/PFC83h9N9JlWGUNsKNHS5rEhBCSv/ecUG8sngaq5PBZUH2cM9SB2aN1hx
J23ifFnXqTp1A69Yv1QKrPMAYfhZ0MPcCYjgUOAcvH6lvCa+j9hy4uXyX4ekZHAfh1ZJrRN4CNij
wvVYzSCM5K2cnaMel+nf4B/q9XedZXpR9RiqzrmOnEdv7399awx36agmnpsHFQcBWUafbvb/Siq9
pTJG5awZleosxbNGKdZXSqtf/TfJG+KuofgxpVwZYUoQzdnPbODqNqIjKzVGRyfbosLrHmpIoOCc
iDMlQ30/3NOE0xyU7Pqi39vK5cBpKJnFARJGI0tyf5wuNIglLcXxB2qec6GBHimbVwIC2o9vJavw
xmcgJNn79E/+Z94UPdm598hUvYR0wA1e0YDUz0PIywJd2VI8wTD3x92QEpV2zHwBaGbM9rmTHf21
kuW4cc8jOxaixy/Y14ZuPFpzSu8swTGD6DGuQ/bmibvZs15HaCkCCezJp2z86iNECx7lXemf1bn0
Jo6cEgvmB8du476nntWOkiNEOxHn183vW0bRyUo2kG4LvgQdbpdGe1VXumtAQhzzOWM82x4Y/wYk
KTeISuwWDEQ98nwKZZnXguYfNBxApjOUm8+6LPOb5N8itpasu4Cy1oNGWLKEdViZS2xmJe2VdMv0
3+Y5xaRXVnhn3wGO/SBZahm5fWIn19xH690AO+POaQj42rs5Sp9gAJkN38DAVuv36hMjew/Q2l27
OhP2tcOEl+SHpgbuT8JbZSWszrFEao3cqeO+ONtXtZmNOVcTeVvdwKf+Ga+MAb7/o/m5Md0eXgNl
S4tvBaBqD+pGwuqXUQvTsHetjEFMS5WBltCo77VnGHA1RGlw0X2svw0Oj6Yox1/Fc73yU1eNN/fv
tdETx2AAd4sTng1FpTwTu8Xn7sVZmQRhackDiODlC6rJm/Ipe1UBL4KlEVcLgPfRyNFfnGoWqiew
CmIQJ5IeyztrlKjMkOJeKXj4vZ56EfQ7N2JzPphPeA+mkYq6RsOy18tHAagkFkukcSjuj163kJkw
ItFpPFTzZKnbLJgUtAJLutI/C9vU/vsVBo7dULp9QXexh7Wm6kOUDcLmJXlFN1op7lNQ6gWlJDTl
6j8sueMSWqZUVpckhfYOxPzNtkmAcXCAGxWBKtV9D9n8Pv2Klihj+tITHZCYqSKUM6TOjiSM4CT8
wYsMYXg28wLEGjkg2bI2llsd/Iod8exGlLMue5vyXbM0Dr6T7lrylimY9l0TzC25alW/RV3FCHc1
FAFdv/zBNr7vv/T5KArPLwk5R+ymBpZ3BRu8Gs+2uzrcWvcsDxSlTKy8rJb3bK8AlWpxwat9uxse
1QBar24pOOLhm1xXioBVCqG9+c4AqI8r12eG87JqfNXwCzXxbwfiIs7SCKJOhLaA3mzPpVrX91hs
gfIsLVIEyMn+ALLvSuIeRjPm+wlt1ncf+Zcp2ZlKzBycjHjUdrQ61iUZxaS1S/a6VWExa2v5r8L0
FMk3sWPVFYMrHjSxjP5+G3vOfWW4+ItzGsPz7B5oL4wIPS+sURcHJAIa3Ip2OckpLvPCxOK2hjFZ
qz6YpZU/MbYk6FUzaXS1SQRIoBvHjGN5AR2Ng6Xkbkns9NylrbhqnEsicoxORtQAc9kVbNH3lNlL
Fv2gd6SRjCkXC1mwLZX089PVsd4+aaeBQzpRk0dHelRn4j2dwvsBS9MCT3yquRkmKCJgwdjt47wO
b857Z1gPtDtgqAYmanlRqW5x/LBrOmtP+HEglsP8c0/APC+lg5mcZIqw4cSGYbraMFNs+LM5oyxH
pCbga0iM1JJ0kbJaiMYQknxU1/xYFt5eBg8+66Kvo7gOPu7Eqtq+mMC6uHj6S4voRJgAxKmU+mw1
UM6u9kDhg3+Pey/d90mZbRApj+/7Cw5TOo6XAFtERKFVZN0LO76xnhDj8d86kvLoMNstynMCECSS
030P9pUvp6zGhBeLTCKQUSfbaQYZrTB4vnBwGET6bI8osthDatLn/w/KKnFEabNp0KpP9q4KeX0q
HhCoEXSV8G0t6b88DxzEsRdjvZJkl8VIJ+Xo/DnUxoVYGe7m4Ezmo0ab9W0bxAbtqE+yHSRg6722
Zx3pjASp5h1vOk7j7Rx+nr5Z/DTW0qFlww0JwSjnIZnMSlzLEyPOf/DBvRW+ZcO4pHGIavHbhQ8H
6TwiGW9XSzSaqom/wmTJA6MHCvmt2tMlO5N4Lan/m016s4AUCI2Fx6Hhy5oZa2KfS0uacThO7erW
xWGj7yvKpHvoG9TSyE38L/w8Lf0boUsmfINfzOrVsEVoB6FsV8HAlFxYiGsUqNAn0GFxvYVKb0yI
5yRL+l7KtjMQKa4RJJ4EyAEsAsEbB9qMFwJ6HNaBunyWSJOgrQkf03D/LvmTjIfJ2idgT1WFXBX/
7SL+35P/zys9zT8OjsI/FIT/PhvmzoKtQ+B1ha4UGINT8ZtVuFxgqR8zYjdIBswSPvjss9yfNE/Z
KsJeYTXIw4EgdaEFuDPUeKl8+er6AiQqP78rmD0FO1kvZ8Uocng55n/Gim+KDMzI/pCh9Fsfw3ck
hx1iydRX311amQlqoK4LAGUYCY/rOMAhgxjDSiYLutIUVgr2vF7QOZ9ZRJB0zWB4pY90emUanR74
ORwMa2VOhkLcy6ECRr9TsBm5TmmV98D7dxsaIPzkGyPdIT/Ct1BRdUPlj1PUnc0V3AY8QIknkdM9
2p2TrxfR98hkNEfyxk/MczUxzRw3flUDEKwadmur1EDuoza/hPoxLvH1+d75A91QP1dTgwHEdwdu
arKNyzSnnb7K0aQAgwdPp2oXNKjzmf3TWVIeoQ9n0Ln5/PIWyBOvQ0SWE4lVLqh3HUpBYB4mw/Lq
oWLaqqt81fqCz4yIPIirMQB9vLsh2O0QV3EadtopvCvXvWlcTPKSFNM4UhLxLnIZe2sbXtZLijXO
SD+YhWor4ru/Ude3+cjLC1EoAPDrvi5bvohRArQqRxJg4nIbE8HTjqnbjB4OKRM+Omo1wfXdd+Wr
tPWirJs7voU2re92OEAAErl7ZNVvIxKQG9yNm+Pr+pnxtd1qHtfNlFRkTnfre58Ilapu2anyXG9Z
1sA5r8uRdVFvDQFx20PqQ+F/Xcs4cCG9YBSOzpWmGVyctmsSE2l0bL9v+2welTr4UhQqAVwEUKx/
L4ZlPHDjGIJRG9szV2+IeYXA57QZjoe0oNCobDkF6OHtIAQfM9sKJ1YQdUGR7AgCtE/xL01eJJHJ
aTmuVw7fqAQtnwASYg7apF+ldPdsor7+1uuJleTFQrb4nH9R+1GX94t8nWELJisJiPZFzqElvAdf
kc9NvNR2BufDA1bHRF/XYLL4Hhv4KDX8q7ukTayXp7ccPj6SE/kL9tp7lfgWxr9wuHum4t9hNqD6
VCXuUHJ/V+6bN5Fbg+Fqw0AkL/G+9UZcyHQud+E/b2mQbk5oCfEFdky6tuT321OsevRzFaK349if
0nGZvXoAYOGljAjnSlC6oVa7R0ohxNNp1I0FfrSD4t60M9hqwofHq35Xh6j1gGWn/Ozd6UV7q7YB
hNUulydP77QHGfF4BF0R2m4AcK84TR4pG1PMARA35AbUzxqftrQtWLokUann/K7pjTlsuykfPSbI
hz4SFbujrNiboZjfaZCUbjGyXunjpIhOlRBolzSL5C2sp3gzGVOanfMCx10ggrHpJNBQxMThcPTV
UpDn0sn805abed5KwnOv+O+BOIIEJh2dcYREly0egaEqK/c1zrn0V7GBu3rRV6ttFva3VDS7ANZS
VoaHI5gjGeV/QHPs0+Y2Fz1F3SFQRqqO7GCf3LGPhEsKINmgDXAbAjOyg6yEoZy11tay7nBnA3ct
0j4ILl45n3+qGz7N7znexoBQn7UY48XQJ1H4BBPudqmeTbzo/KknkM85PqXaaLKaISs7+g/7RtZc
tvUJK7bEJO02rgdAlNs9cyuRfRdIQK9mt0OERv0FZKag6yL4Z3osUsHjbkAXpenhiTc5xSbEa9NV
vutrlNcBi9FMpwVMVUhMaSDRtCdzpFH1GFnALe5EMCc1AE89ZvEPqCXLiCWrOzwjZ4fqy4MYUuyq
V1f1c2GAG9pPhNde5ZERPZA25C0vkg3tQsEHEHVrrDcbOZSfV1dwVWr9VUcYa6XVEgYTpeNx/RNr
HQ/z/4PKhD8yRSethIPjcBdIQEwJbSyXKy+Pr7PkFT9OFKIgPmZJmmheERKt4QS6gmxZ1/gA57KP
QSRETboWngnlvtdAY3VNo77s6LssCnhJ4k1MJM46TCtwVPBv98wS+RGZRq2+IWWxHPvKRyo+sQgD
PMzJalRnt19AzbI/6WjRO9XOiipQ0U6aooziGGqmO+XffxXvWWB42KGmhR6pr7VCQiJZS0UaT2Zz
0+XqWuttxgtoG71QDYE58st3JHQbg5JxfjpWM8km6JemZ7ytodw6gCJO1B4HI+cUPCDnWOMWiqQu
Iq4=
`pragma protect end_protected
