// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
AdwHToWUg+OBXth338mQRyVKhTcI1J1EpggWs98O/ZFRye0btN5EBJv7036ZTy3nUUWKJ+gifnW0
evRfLJVsVtvguF0Wq/XZ/4Preu6/smZo3Jlhf5km4HA4TixlVEO1acGVCWoOxLHxJawe29H5QCTb
fmmsAPNDTqzkhdl24Ukj6qkYexZvF+dxQV8yvxU2WFTOGIugl3elhfLlKGtnWJMw3OpXHWKaNJ2v
yi7vggR2HARjWNVI9Oc4PMr1a6elcK/uvt31XPOssl15asu1UgyTIN+8b87jJNu7TkX0ZttTOFhz
kWkGx05BGr/jGXLOH9I99H9fbQwasDet/yN/kQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
8ljhwUGfrg24Fyyswg4GXgfVPHbSCvuK/OPTEjmc9mjAriWBQCCsdEovpRtA0S2ZYVV+lcF9kO6t
DK4HO4I3OpAQop1gALdCmW0Fcpk3Sc/jVraIHvVf7FohANCUin2h9D1AyHBL027XEaQS+V2V56rY
8VRNJbj61lntBeluzos7B95i0LeKPL5Xxrd+KU6c4RzHS6uo/khrs8ZemJjtxkWlrZ6YnVkt4zWz
cGBmvaNdxkk7izTFsqbQTm7o59FUItectPRpqfiDKPnooJwjZ0APSdgP5MdH12oln+9rR6P9brIg
LT189XDxPAuSyFbiOZt5gzsxcBZg83/VAoPGldklbuFImZ+DG++VGWMlnIWG/KDns//kOcK2yPW0
8YZNfsGnHOZJWfuzF09MaX09gLI8xnldf70i7eY3C3JmVyXVz6z5huNA+aY4/Hu8DwNC6rjpPcGG
jH/9BaFSI7Kd8FRpSrCS03+GPFGgzbsL5gPi39vKze8LTPuE6BzVUuLrqv+KeoFijXw22sjCp1mV
rrVnBwy3iOHDCwv8FKUJvebDpiArPWflY3E1SAb/PcBGQ/JP9B1WM/38mYDeIOUx9omVowJBxhkb
NcXmAtNUA/suLFWyMaSVnZm21yOVwtBhhD6kcsVNf5/YNex4p8JTHUhWE6JNuMdZvQwc5ojqPgFJ
pwq4nrEHnD3KSmO2AvN8lN1zuIocGuo76x2U068A64l6yFRoTtuZ7/syO4NpHsAMnw//7JGS+P5+
uOpayLCl6lDfWJc4kQ+CAQvKTdzbf7poMaL8BvfSrYHBRtipxBzooLBzXuPQ2H+j20ViHIKeFe47
r7OfEINvXb6IPaVvGJelcwuItORkt3jH9r6IXl8mKolIzmUscLLihxxacf8rLjKlLbCvJYO0QlXt
gW7JGLyDmqytlEvQW9pPrNTKgMkQaNuUykquWZ0yoTleuqSVZAmwhaa3EhD0fDrC9NeoYSEP4gPH
1LocxgKxqjdGY2NANi+BsJdAQgluaLahneBqwPhyfJycDuRPfHPthav99ETYRQ0tzoHuX0bNBFyv
3MfRvXipUJpNa0p1H82YqU0d9Br1kt4rxbQGbAer5oGEiCAos9mI17NRxwtZ0uROeZUHuG0rG6U1
vmGweANW6PEaOIiZov0LEitHxBF4/xoCQZopjZl3cBpkkMKT+2zbmxARg4oKSRq2w5cWAm1zGlQH
rTlWo8Lv9xT1s0Jl5oTlLhK/EOjMNY8asKp9djh3iVPK/JfgFAlrvLZ85AMA0c2290UYUaUvdSLT
KWkV4xACzCRNEa7lgmTWsFPYjPbEudJziujtH5tWUqhEH2S+BY0Hxot3Ygclw0A9n/HGu+eQUOvC
OB1DCZHC7yFX4QKW0WUPCYbtKwbzoYsMGt01fIEXEM0Yr0Ya6sFSo/w49FZSrsUJLiUI4wtdDSo0
2I+1KPHu9pFTlRMLfyQwL+7tKDl+mn0sg8DXW9ErK7OjsPhuar6M9kCrpr1i156HOFhQ27L997DF
b1FQZUtxyOY5bI45RWT47DTGhJRynXwTpRVsGSxq8zHt2bmeGRjZ1v81oW41dHG0n22ADx5yUJmX
NM/NaI2OrFnYXhanbNDasuKajr4lisxSxWFYmE90uHz3eupAd659imTJGDH+cc+n3CmurSd9Aej9
45Pl5roIqzNyX+IMzcBMJtLCYMZiGSWHg6dKN3VKdbgNCPppWEWgEUD9o6mIqvVH5XEu/ZZQYOWZ
GacYBPTPi0MkJZyldzo0KKAHaKGOQ2XjBix+OJ1OYHa+hVRN4dmXhkB4KDMuLdixQg+K2jLgGypE
+rE4bOoilOwwmd7jvfOH6Jwb49HXa0DUEqjG/DNQPF2juKFN9dhxDPX1jOvARYcGQPDU1s1+DhP4
TFwCI7QLwNljrEppXCY4Pwnk7TC9ZqzpsrgiriSEpTkPHt8whQKy5yqL9t5mCM5gpbqAkB2SAyYh
GbxfPUyKDuvpSv6wOGJP/TrYfk4PEQ5j0mhcOgZQybFiXL/t8ly0P6ZuInKqbT0KeLs+bkNTqhYj
9GfzwEjbUzgq0+3PtWENB5roibwSi6pGEYOZaGyZFwXvInXhL4WuTM9cgWrCbFcR57j5p/716swT
2QgfuIki3jmcPr+a72liK7Y/1yVsY1Z4zfQj7oj3MfxjLniyh+frszQLoo4ZUBKk/B8uQOeihpeH
iPAMzlAqP24jANiUGIEYfiO3ciYDZE/2vx4JA6eBvqKKpFNVUV02Ghgzw+vadJnG0liMOSubPHj3
MHTnSUy1AAxUPFUsreOOMpgwhxXrfNQpt+2dNLMCwo1pLkr6pT4MKIA1mPXBX7MmOddLjw7eFt1S
8Rp4h8wWr2KTRNgDmV2U61yxVbSi8TqaxjV3YBfdRI/Px3IbhNUKIQ5DzcKid5PwbzBHbz0cfEqU
NSzgaFJveCH8TsjHg2hm3zOd/zD+K2ajcQ8P1gMvqTLaOzQfnqiLRQv27ur03AZKglPScCjsSVpt
xatxbyxB232fIvnjr9uwMcrtpxw4f8MuW0rkkQBP/1E/+LFfz5qhUCJOVRM2u6+kKXM9LXORc7fq
0jqOvcErd0UK0e67OBkLZUTWSxfnJ+vmNfv+6LqLaYkCvDTWZfAaApwZMOxaD2rhSY6RfidyYaUh
c7sNb1CXFiT1e+2qAUtwb+vg2cITUfhbKaXpbfu3GLQu00aikHZhNkEfCxn3eAynzE5CfE13KeWZ
Q7Q4nKrReH/S+0RtbAg/OsqPHoY5Oid9zqLsPKXPGxYha94nQzQd9yhvY/RIRYB+kV0jT8kawnSa
aS76zPonZOpajfntmABoDMfy3lq0jb0wECcAOLgU2ge3ALT19aVSHixwgNu6WYu3CEjfobrQoJhR
nhP59ry9pMGKqV237YHnqC6oq7Pap5+OxJU8jQiZPn3ja6044KigNjdASZoJ2ruJW5xMAab4wVZZ
0gAequ785lHotRBhApdmvyLPsap+hl24m9RoT1xau6aRq0SAbbpVQt48OlazTy5LA8J+glb+Qt3T
3doECY+0rUnneL1iQaL84w0ZNDmzcMHn54P5K8vE2TSna1Cn0cBAZFbNYydHSblgLti+0ylrcSFK
zypjkGTsBn1sUVRlzjno8IUO/fSQctFx8p4NzVM+PnUFU6ChSNyxxZSQWrcb1DmKVKL3OaptmNR5
KPLqUvDtdwAK0kPugmITfuW56EidEDcqLrVWXkBSjdE5fCj21MO4x9IJYD6JGN81TMOVBFJewzx0
C+AIN3tIoRy1/jbcvu/1+de2dzbCmoMPbmiW0mMEA53k3oMx7WK9x74/EwzPU3kY/FIESbhxSR0H
6pyqNiujUwLe02C1P/lcikFeUGA693R0XVtw4lSTuKyl16cAbGhaNFIb8A1MOSc7vRiE+180l+U4
PIZJyzAP+6m1qriniWKufwQ3T55yV57cxENnJdgor11p1GqhJFVRwRm2n8tcIGcsI1m/SDVotyfm
pa2t/Q6UfuZeRSYUydYEmjR3m5SmqW5MxMp4EDh1G/4zpbYe/yHGbp8z3NdYfn1xkFwOrKU/bifQ
9FeZ8F2BNH7Cl2HzpYB1Z4lZkHBY+FsbAyy7BfXKrGUmM2gAy1AvJgtbEc6s1vWv+3Ot5fpTpznr
c3VOUofAkGtN77Qv2h/i4iTpcy+Aakc1xhblXha9/c/kHA6m1vgWlJ/0utnWN+3xR5liTkj8t+AD
ZvU2C8hrElIw5RwANw1ipI7D6MVi6Bczo5f/ZQ9MrvmzoNyXXKx6I1y8haEZ95VbaSUOT/Ry+j5v
lT7eBEuHC3De6UVj/85sfHQUm7uVW2bvacG7PfNdf6x0n4hWbV23gL5yiFwPkb4lwu5LFbpKqWqH
DLI/mG9tLsy+STGMIJM52tVUDhVdQdmWqnvazqxofDt2JLaw6CQ4fGCqfDoAAiv7aZqVaoy69P9W
CbuPxXtwNOxr79S4uwjoEcF8zH9jYmjqCosuY0EwOM88oIn2vT2i4wUh6NIp5abYH/C1pl9C6IK4
5y0qRldUgNeHvfAhgyAeSrl3BYfhmFMTsasRSiYzUqzbPXfM2q5EHJDaVb4JNb1+Czr1pxzE+s/f
CoohnazcKBVi6cQESmJsCEnkPTLt01U4GAHsFAdI3Uvq38ujY9FVwr0mf1FPdvfDoTiXpsbdATOV
BIeVQlaAw5cG72L0cKld7efcq0zVtL0OLdiDCdbrTUfjn7N/c/Nolp19bSTJnoU9kfrMLKq5GagT
Jm57/2Y3dlWvyGlHGOJTYulltsTHiR0X/v27i6MHREEyFtWwMJBElldY76DI0wOP/vEKy8dyr9uz
Z4eTGC2CAH6jhJlfYuEPHngokWYikjEnLwR3NqGqg4rKfuUBo+tbvvQyRERwA/h0QTTmBJwpLsab
q+sR9wZA1RJwezRkAaL7xXiZIzNcxiQWdBRgJaR1T++rQk3Q4NtrZ4HuXeZvT84/bpWgUW64tekm
qIv4rY9AbYOspwoWcZxbj4CiTniIxGmTtu+Yeb1BB1cMQ7sCmFGXx1krmmb3Ijb4Yttx8CysouI+
Sc2gYCbY9jzFVLv63fQs6/AyAoc5Dkh8ALMplVO5gZPX6O8SAlyDO59yewTG7lIGKo/dWYgTPhF8
fpjXMqaEiZR+iyA+gCOJkU4Z54pFP6+t0jrZMXjyijkeGHxU56NpaRrNuoeccjRDJPX/Jw0bAM0t
TSRe13rFFfS7yvb8JZ7r3cZmEIq6mgXmVIPnVBlaXb7algojhNxbiI24S49yCAwbl9OCXqJzlvFp
5lwbE6cWoJmEUrrjYprSOO/krbjYxvoZ2l4sx3nAaO0SZzfaVaUdjMZR9DMcrHWVyXPIdZ1Q16U8
sjiDIx9chdjTe7BR+kvjtHMO9y8u8ZxF3T3Eff1br/nYd4XUDGdp4r6GbHn6b8hR0pbJ28TJEkCZ
E7H2yuBZYZWGTH51TQmS+X3LITmRcKypwatmLzKDYTH8PVsDzRJNyZIWfqepraLexAv85yhzETTz
qqmI97Z2H3l/OzLPz4E53EwXxSa38OZbco8UBW+b0AR2UfHksR6lEfPj1VaCkUCpd9OrV2h6eaKj
8Djh1pV9r+76PpmnwShJAcyC/SBh76iN/I8l1Sb+Cc6KSroKtI4EgncFtawJ7RAIPJWYY9DVvQeD
PV7GB2tAildkccyhbNrF1HK0A9v4236D8o02Oy8Ub+A0A8Xm734VlBnwRD90xWjCjTOoX8ySV9S1
k6lR/UOR+bDx7ePI0P8O9tUOo+Y94f9kJXWReR0oGMqdevBO3lfg1la/lNNb5KA6ez17EPBqe1cJ
AD60AAQnCsl8+ATaBgDqI9STHir8LX3IRu58Kxckti//wpW1KRiFSzIW+Fn7g0JmUhssFldi57ZA
7t8O/t3FoTm7W/x5g5wC2eZX/QkiAO0uI+ahh44JDsn2x9fjgx69q/zEOQxltwUYun66zVUuBPPC
XZh0lpTu6hgfXksb/hD16L0AvBnp5xKZViMz+3X4wXFqnBOEqTrN0DSgr6uuSm1qSf3qK9gg8jIX
j6DcNZ58tNNW70226prA6TUGidKDzGi6oP1twCJ1xp979NGPyhEB4mMd1tfkKg+2jDKG7gbeov0U
bHJeugUEoBXQZJVOI1QvizuMUlpJoQPp/Q2gBOm+Froi5+WRwxnzennT/jR8b/Woi33+FKSjt20B
tjfiJejuOB86iXal6wbVhKdJcWwFbxsagybJ0YmpqzWjpH05qESqUoJPCKZVBO6n+qiO+3gqld8n
FTISduNAWg7jFPceFpDOXtowZL7RafHJ6vY7nntBh7Y4fC0jsgH1QHogdHBFgFyf7I4XyW70ZFdo
D2RhnXr0E43hac0KjASOT9hWOf+npsA1xR3Rp1wg7W6Vp5IH3J1fAL8HxoA91nVGl2iT/p9Jy0ni
1oOiA3sKEXE/LwI36j1btJG4nTdIvoGsq55J8h6CWbP5sXvAAvF7BMBPYLBXJFxgS14eii70t1ml
cBIZBsVosWcx/0g9WjZRspt++lDgRMZlnbTxCri2RhQnSd/a5qwQs1wWEWQmKf1gJJRfWnqQD/dm
3vV8+J+TTZz8TYgl7zD5rKm/nTWW6EcfPOifgU/6Jng90m7TsWrH7VhmNG0yVx7MXbsYJiPjBc6N
C/egY3pc1rjLZZDOs5ssDC4KmWrMsRwnab00atDgfZM2v4e9TMM2cwwd3rZaO70CL7QKFQwzWMIO
QwfKSnuLe1YkgzhXI+JqfezTMiWBQRkLXxEzh55m3xKbtZIpGi8qb2REEaXANJ5ZnZvl94nlwbOY
eibZfZac2SlcwPYjVjSqF9ivRos/8Pg9PivaPwxhMxEyzQWoOcQL7mX7EIqJ/j08BqpHUrhPhhHy
2KeTMEKPyBLdPJRmoe5hXlzzS35uh2fWu3iqUuprYHmhD1MB1CbzmpYfoLXFQBJYSi7Lr+n6fqVt
SXQWZ5ye5uwFx3DaY0lNkdANZar5sUnKW5M+0Vby9TdrrefJUePTMcM/t8lvmdfuwpn6myXF7iiH
w0NBURYL+PW5LG+OdVKIlFcPFH+TsAc4VLBZUYqs0PirdsFJSVf4OgEXNQT7dtrSjIUEPKDyy10L
3wtH9Nl8CTn5R2aYdZsnV+yEML3dz+Mz9e04gHiHnhdCKrgsmhEujzLicgl9Qm06JJ2V9RpxT6GZ
thzdHwF57OKuqd5itK/uVox9Mc3R/1HiJtkG9sTuHX4AGTn0wvyqJ0fDLDz1HUUwiCRDewllNZcp
Eq+xmcu3AcYczWup2hkSMEQIIc0afsIexWFMFb+VBNlU2OBO1NMD/LTP1XKBRJ4+Xo2dWS38HEGY
ig8XNqRZrFIMPxMvtJXqn3/Xzug05/1/Uq9Mk4UwEMyvJsr1E7G4fJ0944U9fDtYz6XXjAPGX1Xz
5Nh0R8NhdnvlBKYz4CpsiQV5M2MXk3WQKPb2OYDjyl7TFgA9GzVvy+bqScrBSAT19WIGo2h11yc2
IRaeMsxSSFh4UT43CGMFzNJHQIPA08+1FH7AdyRYBnfZwa2dghwsD5NV9DFNLCeIZZShiOmkKken
oaeRuueYBQ+FDHYAkwz9coZBrTWQVzhyt+wwpOehQjypg1XPMFAIN9l1MHJ897XO2Vupe9NUKBbX
TUVVnxGQ5CqUrttwCI/pG3tFJueoPO2Zo935u44OL9OKrx6DmL/h4D08vlw1XqUk/scq4umtEcrY
Hzv2lfKPM37Q9CKsWC69U/UuAJXXeTAdsatL+ymLCmEnn7khF/25Iss3CCHcOPd3G3jO6+LvSbfc
K1GQ9ObuH6Q9BihQufjyruvmLf8LjClrPgCFInbwO5m9NCLUGHhlizJLcX3Vv4LEXYGrdfZcVIK0
BJXTfcab5mqkbDF93cWQlF1hJPLP6W8kNUtn/nXoZRNWAWk7aj6/q9Xzfk0+xHyIL2l+yaMOMC54
YtY4nVryrLLO+f/DvfPx1lpHPAbftnM2nzDSIgMDvsTJLJL+J2V/scwLYc9nbShHGAxCrqn1ynxv
6KR3t63wlWGxuDlw1L6kyVI6CauIFaKZIYMci9dlUysDjttAud8+JLc1Kzc2RGI4HcnjwV+XYRHl
YmPGikLSgVEqQuKwu8EPnR4OTvJ5vFh+hj7kopr9/S1koJ0fhQE1rdo+9tLajduBNlhl4acGIJgM
2CPvU+p8AQieERMb11Wkduq/9zNUB/rlrvmiTk1FViQJ5bhD8jWqO2M1iIL3dtDklMYsmflW3pzg
Gle5AsPnbYhKjwFhyQ6KSi2wv5CR1seNBXYpOhxsffJ51Bjx0HjxbeIJ66d9wmfs6tE/lsh1tOQc
KViHFXKNBWezGp/URx7sfrQRV81bYGftcuIWrW/e3ZTqNEKnAgq64xvrPfxutB2+EjNyOAmuiMiu
5KO6Ozcixfj9dAf4Kg8cs1qAJ/bY1EI8nCU5WDXKS6zCA0wvp8I7yvajXWdPJTTNQfjkKkV1bK+V
/indDfgf/qTqRh+vLX6qRwB3tJV91lyFoGy/l0F903sLxWbwvaiJ7y1jOjrvXG6o6RpbDkWuWnuF
Wyp18O+Ev9x434dD3X9Iv9wClBFQSNU162oA62apexeiTFhAHWpAshRiByzXqIXhgGW9rnKPD+/0
rGd9oGdFSSmvscqYOrEOYUHyNsKAqEUHyyC9lBbeEh7rJZDY5b6NYSojM/NkMZhE8t8mywX1Aqn2
RIRPEnWX601xHm6OP1wB7MCOPNN4ocbT5AZnGf4TthGZfqSyiI2sLQC+fdpY48Y2SE1PFITeTXwS
UzAFEajpTZppHBCiBHBX+meV2KtdQp7ws6aO/hxoO/GT2y1gkJbg4ospPq7nq7+VyWECmGQIjzxe
h849o4C1up6XSCxMplDJcfgj4RPOvoFSu0haueqZmEquv6uvlI2SO4TwPbrsH69Ye47D92BOzFbf
xv4cfIWHViJp5n9yEoltj9f0TBKOFVD0Xzwm3tR2sr6yiKbsqRXC2V3U89NeeRYT/Kio9oVQoTM2
g41RzkP+nPpw3K1SB+wR3rxkBvbxrEwlCJiiYoHr5X+HSxOaZFBsKWIorK7RZSxaDzG4zgfFVzg8
Uu64BMTVbLbs4B8jg501hWi3hwMWKPAClRrPSBEWLZqZGpDXj/S/ABHMNkJkUlcF/Eo4rcbvxXj0
B/NVJhbfFUfIzXsxQG30NrfGdivxvvM6tu/TAm9vUFCNrjJVuPg3YZjGnKp+HUm2+zpTT8lcxUkY
cmt9KLxR+oUYmQBNZ/D2hdgyhsAQioQmsgx9A+SZE2KmP0IT4l3eoLqIN3NhsPWTDGrsdH63pQqO
rELgR0wkvcFZexp+1BoZ8iLKYcanT9Gy4joLgHSBeZqJMIvXzeZMBgqYZOzvOhFZEzPUsxRwqR3m
T1Tr5XXrjKV39qjpCTqj0zY0+Ta5RQdoxE3MZNwlVxx8yiJZ080+kg1cyruHSAGz5+L6qG1NG1Dk
FXsfbx8yDOqOZHH7W36nRBzNOV33IIPOzlG1ucZ5VEufHdqkiwPuS80zAgLoMF3hI1nwIYo0CAFC
JPkYPSb4rd7FJytiSYDFfQ+EGpd9tnMxsD83Pj5gK6Eic/6ztTqLLuNKh79lqcb0M0DwUXIs2+6J
y6oBkCC+F9+1aLE+y+XbHbhg42e6Gr7Cg45q1NnWalIwtDUfdTfBCdWSjK4fYiDv/I7gCMA64SOm
mMopyscjqaNcfM7JgYU2z8EeZtnqosaX/ctl/XdixjtUje6IUm8L9MCGbbum1KlcbTJntcqj3+/V
rs67QvLBYsEI3ai3suWthucTJZj+GXRjJKGA3z+/1gd0YoHQ7Y2jw3LBu0Dj5msBAsJ/Rs1lAtWD
yYbMAoygXeyATejHp+wAeeUTPWvNVEINXAYPyeYXyKMvc81JfQ3hIM99+3jJQ77OfVZerCw5RZbq
/+dWrF6mcsI7cH4U0hfP5OKA3wj2nP8dgT3aGhZ5OavHxNWtYfDZiA7x5xpkOet19ffF4SqqKZ9w
AoSbm0x03WJHPuzCDisjgrVDCT9lAK4BMXB95I6amyqpoPQSSA9EIDRd3nwuUQkoNpfvYmN/c9Y0
ZnuIS/Z+xsVyQ09jmiUep8KtwC183tBLjFrK2WieSqF3aM+m0iYU6TL8g1+mM2lR/Vo/hEBqM3jy
d32F9jJxK+s2b4LDLDEcoFuuvFJgdaVCLEDHeQkgPM6ucgtJivztyj3N8/s3FmgK2w3mCxUeF9ko
3+GFdbB2+3h3W5pWJ6oHEWkKi0SXCL5VjxYaIgLvL863x4dgDnhKiDUanLY2jSf9HVCET3WF9xpe
XsjPvZTY8XMgIx+o89GLsTpKt2s3xypjzSnU4QZlnFNOt+2WXZ+SI21HA+wksVFoZYtEAO4yt5cG
DcLVoZrIYwSg0VeEvb6PL4jHnXJjeHUNwHWYkzcBf3z337MTp8zuV96/hctHMAeIqqDYnVvGx9A/
ZsQo4BanaiISiNtyhmwgVTlyHHJx6jNzBw09sbxYmgowK5dI6V+O05oIZC/yMrXC2LBJsIpis1Oo
KFkr08+huMfITTyEeemwrzw6aItf2kpItOETtNYGeSUZKRjwyfXLZ2nq7zUCf66E+An6Bluu1BW5
u9mpBDDSzwOWKs9WO4cw4UqFMMMdtk6RZxuVvmahxvMFtVPp6woRFzt2IO/cmPCvuF3ZH0Aynnp5
ezeiLUrccXbF8MyiqQRQp+2/k6zgTB516fackDJeEHmBQTgBuVTzW+Rdjkor/R1eMalEcEEgRI6c
oYFULXhGgjekKfEovvNtf0dd86v7Zl+9du4Cre9eexpWmzFSpz3oKc5eMiQ+0JthrlkRVONSGtt/
3iWJaoC26QK7sLpM6XWQc35LNcPhYDZhDFrPQPjTQpgJj3bJSyI4ErQZ4pm3acwADDp203ELpue1
3iwe4/DXojRoE9DK02rj2O9i1+qf1M6giYlz/+T500qN1xrzBol+DikjE4QdVQEsi0Fl6KbbOs7K
0ni2hyuQmFVqtbpNpfJdom5150OS2rdMOM9X5KFUJzJqM+zhvBibPWad+HTdL5a5FRebU9ohhP0M
72JFlB36941cH4piua9d2zRRA01RHI1x0iCBg9XnjZ/0K9226ZSyXLiHPKITLk7GiIO4hRVgX78G
pSuwRuYzMSL7pLmj6HhWk7H7DbOg3ef8DWtTNCpv3cF5eAyCYmKhf1BMpKy3abzg/a8UvonlMjt/
epq18t9GL+Y5hmhvQw7zcYuZPc8AeR72gLfEf/oQmI2cPp4g3E1y6AtDtXIdj8wXShEFfNGNws4H
PX8sddqiBNu3oBdLnDlBDRrlnpCksTBPkIfrE7fAwdwcF+mNRPRIturiF2uYHWyHx7K4R19ouIib
RlObKuPVYiAthGXG0Ql5P4jgni35+cifmFJqzYBzsL7cCw9EzGQ0xc/l0FICU+LE5VbvkXtkMRYx
pqNsdm1qa5u4kVB14wrw3bfpoSBDZ99J2mIKg7bpAmlps4Wi5pHHKFz42VJKYW87qC7yLp2tZzpM
ODkRBGL2Y0WDa83Qd3bHps8aNFmkYIU0ZWYHKa3iyiIg2HBTnU0YLYlD7jSD9FyrL+UeSFpJ69NJ
smfz3IhZgBm7XzfaBhX8bAj5RXTzSwOP6vD6XVfdh2KYuwvDPoxviy4Wb1n45FLc3sNNySuOxCD6
tN2iax6yKYJc161PH42mmN2LNdbXQuNGyklkMT/pOInyc/TM4KwdcQYDXI+QhGeZmf42gR06ELru
P+RCbT7pG5TqL6djzXHFStFGoirPpc1Hr75eI4mpqpcCN4lS/khEQzXq0zjo/rdsyjcP5r/1a42D
JowGEggJK7/CzcexSnlB18bCFvisFXj8lpM1c8tQanBfIN5qBm1sYgSuEenigV6h5A/BqMpAXbNX
dDkJ+9Sk8WTTt9ZF0AjlCHxgx7SFra4Xj9Iw8Okr1EXjmmup8mo6cOFU8Grim7LhN2ohFnQpV6tH
ugB9yKQgscxEAU4f5vZz1HY8XM6UAFzT/E8Nkh48tpDVD6+8+dB9Dg6f2c6trz7cFmSZnVrJGBES
b41nfN4c1cffsNs+Zc0LiZhTbf1UnJrXokUvXeyHCOo73exet9aP8STPPp+32nGzwugqO2+Osvly
CVECz98OC/MUO0hv7iu5c8c+idHVPZm1A/gibj0w+XtlSklMD7Jdecz7DWhl6mEY9rewG0/3uvMY
RfwOMVHOozKBHAz0SMjhNFzfi6ygzMxml+m+3WXRkuxlP/V4G5usRZkbffLFULhIqvC3wkUdGRZ+
PKgdJnusqHII5t/Lfldo+CfZWEjdthgbC3nRWVnOALSGQjn0Y0gPnZdwSGatD10Q5WlycRR9Axlg
o1IbSBFJRkB5GVd0PPi1fdYvk3XfsD0/LJ1WZatCDaZjPSgkjmNBsm+Ta8s5VsopN670Y2jRQ+m0
83tIYCF1Z7ZAV9XXZ8ru38l8rtFfHJB+ZZEJaZjpVUlOZtPLfjwJMSBVdW6HOvlADVzJytIUAc7i
BWbyyLGNarrBlZ4g0E8mBLOJOX8NnI5yGi9qNWrkwYBJLztQvQiV+Mxc/UIiM2yJo1BCt/53pLRz
W4HvHDI4RcHEAbcnt30GUkv+ev5XtN51PpOv2d/nZro1sOYol5BGjPSj8vluu3atvPFKdUfrJrJ/
pQrCR11I6ks0hKym76AB7rbXzeGJVCQBsIdEhNY+DuMoU9XgniwcPvhF6yFWpgebOnvu3nBfRiOZ
syQeNvVnaNc1VwRi2Wl8r5J7gFm9xuAmt+Yo56LXX5qIzNiV/vR/yGVh00iwe3+djwo2P38JiXIL
tAUf4Zu8LHHPiHrEAXIsaNykXpi6rZfUMGDvhxcPYKzVWRPabxZ1LeHeTsZ/GeT54lH6VJ3F5ygw
m7V0ENr/9fFHsEfjI0RFlRtBVyeOp7ArdL1o0cNgifAL56nNhFNjYjKoIfsOOv2Bd4U3dxuGjpKZ
0CE2tu6qX9IlvFCqS0dqFRPBNaxEhVfyyjG/Ox3K5a1PxPfBrHw2tdN59ISgd6WqEuHSz6Y7ulc+
sslZHe94UjGoiSfZa0qPlmO8XeQlx3Iq7FUBenw14skepbt4fcfVdRicTWiWi/lwKlzzV9kavOOG
zxV5WjADB1ltPJrK6dzj3zza6vpzJjwyosC7ayAEPJDv/witKGnoQVaTdOIvCqX8SWncjn9RMvDm
T6vSxZBVmjKhQOvIgV1F9dZ2twa99rTxbHpGpcLzkqvjhN8mjoSwwKTrVe3bSIjbP01GvrCs4Y12
XQgOKj3CtBNwg3CqxzGpm7FU/838NdoxhcrVYBibZ+BEFpfQWSob8p/lOvOk0gPabQTThN82QTNU
/xN7Ue/UaKWe1wMIgUHk+qw9B3WZBCivHcKZ00g//6kmDp0Bc/EWOrcpCOgM7rNG7/e2k8MUvcWE
wlbXSdC4YoUrYmXCW0sEgEeGajxzkmQd37rOLG0Lyt547IpqC7kGUt5CqqD1/0aed7ofR3KdrnUw
mxHDnan+DpqUo4Ns69WePTxgw6XrVgPH9I5sOzbb5iG/D7o8L8vpqHv9CAOayYWY3PbAXXTlEFLj
dXl1AFzQqgHg/kSJl7l8Mk3FbFN4hUH9q6Esc6NW/NO+2mbH5YVEuJt8GCy06eKj0b9oFQNNJoQz
5jtCkhRf0Cdd3wUrCg/BZtUz6FhxHbiS1d8RSrHezTA6sjzYi8L022fPW5EzVfa2Xbs+mWAK9n4u
/SqXPz0qQjck5S0KqbMeL5olxeexyYfl94oyxwNtptoakQhx5RNvIxvZwqLZcPzNSMACRvZzwBM2
6B41LaHlCDdw9E0wH/FytBcKcdWhkE+LqbTzbKLPZtUVhrjU7mm6qCn8i1Ej6zQPwJahx6a4NLra
/dlViPy5nP6Ob64T6tBhJ5WOSUAQIZrw4lQ8v7gqrjupylt5RmGaxxbRxzAal93BBHpVhdEaQO82
E89D9dJXek21pBibh5qTHBGu3AKiK/mqNTf7bLWydnPyydu6VBNHRX5EgInnCEgOFXw80NdUAmCi
zz1E7+z+U4BBDZzJxMjo7gIz0+JvOf7yn6St5b126ISx1PD18Prc98VYD72xfgJaYEe40MaPRwtS
YOxQQ5JlQ9byw8yGX+22phCtKFLDLMVKfFyjC1iRoN6sATnpk4Dcl6vTnB98fYTJi44YpMF49gVg
zS4fMltWDowJlaT5UVtWU2gav/QsBO6Rh5UZUzrlXlSdfKJqToqIyVz4JKMC2GS0NINQ4iy4bfPL
i3it4UiufcN+UM46GUiw932KHEge9e2GLlSr09Ie/H7z65TMkPUEQCz0VoUPOdnAILkkkLnzmubZ
4YNFq9z5SaxcNVcYnKZYmGmPSzenBECjGa1angHYuVx6wl4aZrljgLWlo9g/SeUS4vm2QCeZQtrj
hVQni0OHlJEdqAF02x4toGNk80fzm4bUx92zg+u2c9xnQaAYY3Vuibji7L/EdAv7wFxpj7t5SVig
iv3HV2LJtbNg+duk3YVOihDTVqPKp3+37AHj5McmNkG/0TMWva8wKxiVaPLxaBNNTFB2G01HO4Pu
t85box7ueCA/59inPe9eW/s+zTl/L94DW5Ba/y068CehT+BFDenG/HK43H4gR40bIBecejZ4ngtP
RraaUKbVRtpNsp5mqiy0xkcbz5ZxrNwl0VuwHhjikNV5QVVTCbgCSk8M0p9IdEnach9kWghoOuo9
aKcx16L5XWZOSQKL8P9mVahKKlgB8vm911GBLa0p7GuT60ml246pnASDnmmDJZWfBQcjzLqtUdIF
OulVE2wFltAOwmPPZ22hJM5fOEcEtkQIp7EsEHg4LEhbvc+L6sWECLCfnMhnuFQJ1nI4ZO+Ns74v
MmE9vR11Ja5zHrQeBoLGxPUowdruFQILALunI8/TSek+dWb85wiieoLrMzBaZ+yfR7yNrqqzgrZh
xwCyPM4UeZlIcladzPsL24duNR9h4u4zRoMh0TcMbNWDHHBtd9JKtn7ACWyCjmoxlw9861GpNaIc
zbmcZXlTGbkw0o8lE4bi7zI1Vtx+kG34Cus5Tym2xO2kB62b4WUc7qCC+CbrXTubbfwP7URPMl8r
/7vw27wXgcMYITcXVyI7zw815rGbbdBwIWjCH/fKF8wJy5OgyzGx+e6l1Th4oK9CUyjGxmyaNXPW
WzSMjtvrgM24wVkLZdbDBnHHjaL645o+59OhdcYUcP0mxo3nkTs4X77Nvz0q1R56ga6rfpYX5QXf
OTO5uIyao+pzf9Awy1JRlPWdN9trtVIafZGEnDruTSM+PMmbtyb+k36ZFbB4NXX/RQWJD9IIT73t
tgRPT9FWWBV4axiFDbVBF29fOJqw6l5m+qneSqavWWyrlTxZA/fg5Q+eWuxj92hJQnOnfdid3L//
7f5zEbRKSOHPIuVMikmzpUvOJbGumO0OTip9O9xiIxC0H1wwKMbWcKKpSGENiPEdKeWNltI78kqz
EZNwxTy5OxTwXaOjHr5zlFRHQVsGvQfvsDAIotdJBzoWgTxgkSyX16o4BKZxzNwRyPhcaNlxiTG4
gpfB/R7GYzWuwiBvbdFiv/qfsXiCyT3w7o960eQvULk4CNZWqaOXy7AeOikPywVuI4o5Tne8vvoW
DrYiCBOLPE/6vJh7MisXjoni9eGqoTTmJ7aQMRiFp+JJiNlhBiYUHyb+VDjdLF+wbCTnEiL2paSG
Ml2x5qkZaImJQdNjAbhtvmo8iegmZrNAG9BxLh8kFjY/EMPhTpA5RBWKLPYsLl0DsynBqIdLZ1jO
hbel6hEbYK6yl7SQv9gSpp/UoLr+4nd8GCJBfmMK5DBYR/B4uST0q5B2s3KuW8V2QyxlNzO/35G/
4f7OQi+sbzhVHDSor5u05kIL/f1/Wv0SPLHkuGiA//hhVP2KWvUn1JE2FH0l2o38SUbnOIDsxkto
rAM6Uu4w3GTZSZ4O+b8VMy4DV+0ppN55jA7IG4JXosTIwiqxEKNLtPALSCoaC43za3k0mb6BQYD3
vpQZk1/y3G+RGY+U5hSAVJIPdn3iobtExED3Clbu/IhIyV+8vj/pOUmexkdDI1Vlg16DtsSRy8zP
amw7FX0MTZAZWcLcV1M6g0NqJSGxCmnZ629p/0ccEMtVX58TPCeYgywN14uh9GjuM3Oc6yh9dZCR
FAUfDS8r2Txz/UwBMMY4+3WYKtCN6iaDyQjd5idlWTiMB79o+0woRXO2Vj03JCgSEApfcLCUcaso
WzJmWmo7Y2fYgwD3RjRru41jU/UnPNfQhwHxyc0e2qBYMBCBMCiHQzFeS5LQhaFmOxIv2Yyc+dvp
1rK46VkJMfx3nksHoFeGGXWvcOPAHOX9+7+/3gnh1aQdkCqXPKh8qGrqfuS4l2hSYN+gfchUyNaL
oUCi6eu1SJy0jUMDd+jYiO9H1xLkOlsbZWC5Frt3Z2QsVoUtli+EjP05u7gR27tMJujBMxdVAaxH
nNhi/nxaZ4jMgotOhZWFXcYmAD8mMgJ3joRTu9vduD81KoIOcl/M07oAF7D3DaUqUJ61AlfMy08e
XIlX3r40R181F1ZXq0MYpdSOlaWvJYc+PyH5hH3mVCI1lIqnVRLsSyCYWkYx89op5N5033TzVmnM
C71Nol1m9hLDhJZs2/NWn0yD3qDJi6BDLSw4rQfgv+IMjiNR0AQqdEMqUnVIwNZKSpZs6n5zkTFE
tUjvgiDFMykZIu1rwrokmNsWoKQDOERa36oMmzUyewNiiBgKY/pV5Q1X192WbAodpbzfvAzeWRR4
dyIU4MwY7Rqjb8374HbbCXlj+0Dg5BgiUTgQFURqa42uW5+QGm1AUqPGnvZ+xRxGaY/VhB6wYEvP
hf9VkfRAkYs2iCc2MuXi2shm++ioFOElwN7EKKOyXbHInEW0bmmI1iCgREJyZtkjW+Xckw2UtksU
n/cYiHif+lP7R0z4qoUet1TXtGtJYJ/l7pWe4i4JPARWIhYRWz//nQOuFFJHYlDlA4PzzMlr2AYV
qaFN7WrcN8rbc1Pw4gYsKHD2tIjfSgu9tCEXRrg4YSACdcfXEp6ARo5UETI50gntF3QaATG7OMfn
gM9MIDjk1QVgRlJ6uvW8AKNl5b852njosqyLV49zkGZBRhXE7IU=
`pragma protect end_protected
