// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:01 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mg9nMnpK2Fr7643aY4IPUruPnu8KR9AF4XL6ruc7dPsTS6VWyaak9NBVK41j2G1J
yvZGyZOgpxuOMYMnn0GIoAzGYqDckGJiGupfIdX+/YAb2e4BM3Jw2VF71KRyTeME
qNPkNagj5HSOk2W+uepvoQ+wAB/uSQjWE3He3/MqfCg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21840)
vwqqX+vDTsrTAUz7IYZ10/+cZSURr9ee7DudNJcp13a94BY9OVRs1fWs29x6TIc7
62f4bR0XR37whFNNBjX0kbbAq3m384F4atmextGbothhRftNGdkar5cmUxxrQ5H6
cN5bfAZBtazozS+hFb662LlnRvLltCivRlAWcZyFVZwxws+sPOxHlAyvS0yESIUk
oxSwQPqVpH9T2InPxIpcuwXcO50X2+ALFvgTjRKluK5RS4yzsxlk1/ojnD1r5Uwt
QNc4V5ihk0Z0zR2C67zNkEMn4ehKtMtVf75pNlj1DEKwqfw+e+a7REX6DlAkpl/5
Q0JRO+AQleEI4o3AV3ZQ2MUEQEDpBrSfbpL0+j4i34TtDvbJl9CdGCp4/x7IcSJ8
QukifEIaTRipBug56R4B0ym2ph+Xu9bBp3eyppkZvEZAY0JW0Q6ZhaaKCbpZ8vkD
rT89++Wtl6CXRj8bQG/b+PheNLvPxKP/gYFPEKwG12JUiCWQ1fk32CgWfmBP2uEX
rbzzCgz8adukKJMXaEpBE62EQ4mwnXqXSdvVFjZnhECvk5YQGJ6zm2sE02cDbWF1
6yQk4usdEwEGjys5Duojm/RM4h26T9hjGokcgdU8fJ2FzYdCng5aqcPvK7/ts0VN
i7/8QQMLjFt9cbhyTppb0gMpyIqWJbmq/cw6FNBPymLH1SZ/+F/9rR3yeX5FlnDI
XZAKS6vf+MJrV+iFG1DnjmLD5et1efl4vPSLqv5UISOOtSm7Zy7sfahN/KwM1lMV
HLnGJsz3A1mXa9q1XLiHulclBAyBqX5+OJLdLjQ/KvjRPi9ofPZLUAe8MvVn40xO
VnL0gAqrmB5N/OPpacomGzeXUQCoeZ/0VYEdQLP1hP7P8qFnYur8A1QDL/FN+Zrj
FY1mKE3FKYpTMt5/27vjhgzxhvLitLngdU08sbQITCijV9KiW/tDuJ01Tlsafm4M
5n9QueXxovRTeLZJIXLWe48xEoTDn12t4R4dWgfTHAl5zVY3G+h1tRR5fODsAAzD
EOw+JeL9QGSb6+/fe1g6D5wKW5Ulo5gVMFH4wiGT6hpwPQq487pVm5p119sPQYvS
oI6d55GXp542I1jD3ho73bftp2ZlEwJrQhwZG1C/h2j+AHr7BLExNAMwk13K5ogi
5doaauT8Ew+OBGyA824gn5X90KMpgtAHtzM7gl0SYBBAd2ev9c85HaTQnNdoC5Mb
opNhlCbVwACCHfWagT97qpRHLlVHztGYrbF2JnV8pecd5EIRuqGeTiySCydMHSUk
8M0ZblVAdEM1ZAQbPGxoV8Hq89dC6krU737C8CChkzuWOVIHnlruOd0Qm6dSXPJL
gvC7phc9Qjfmr23yc34BdE2k/CCE+ITQ7fJAMkoQW94KSiRaUKLXRaDONfKqpR3M
cbwk4g+fSdDhyQQAI7zFsSxWdbiBDTUJQJ1kIMtQaQplO6a6NtNQFXhmhIEKZ5LO
j1vGVSKcEMlLL/8p3pEOh8XwpwmjPQ/dKK8SY89DnX5SosxKApbBmEgPRBTbb61m
h7pVROSxYugavzbyIn/hQ0J682K7VHqPUi4CtAIy75Q0TgLxXi4fBgjnTRqTrEl/
mofDaWLAgdIsme8hh5H1fd8ECjpxea11gkfKSRmDbGEshq9098GzkFi0jzeyeqG4
SMAgwf9TTCGlANK3cLOFgwvW6Dy5lmHFHTtTKIFOE+SyEhYamKX54ZYRlD/4QwjP
yi2gn5lGHjk2DNIQ7Q71iB0q7Xv9IB7A8yQLMJXhobpDV/RSbd97XP475PFLajah
iS0Qzr+lJK8JuStCiyBNWmFitLsoq2N3RbfGDxINhy58xWpZjFNvfQEMCRQimSq/
bCLT06W66sqF+2Lzq+jtjETnMO4LuVrssNmPAy24ZM+56oV6LPs/VYVq1JUG1BpE
8v5GjntYaW52tmv3aHRlzSZaScSYEzCVnMvfi3nBzxw6LPIJ8sR0OumWKcLh/bs0
n8Ai1/GBvcivF0ypirWokItwXbVm3CUk5RFOtvbjLWckt2HUp/6SHk16qTX0OxHV
EUn/X0nl3VyhZ0qPRPVrJR4yf68XFhQjlV7W3fss6iFtn8KuDCigpjSUvdRrJrf4
t1HgEpTsb7HugrwL2v1tige7Iir2INjGzgYazuFMVFVvlBTIRM9mCFS9be5NUgmo
PLtErGzp0dSSC0er9slZ6ahnpSQMjRlw3JHVh2Xv8Ee4sTFgTlHP1qe2XvDHPBzb
cAGUTTWuDtKJTOjjHV3fBcDXNajkT4zgakmGl731no1YiBtZfm6H2ZNh8RxXhX+h
HKi1OzQn6EN4Uv+p7JoS6WnraNAyBPKni94UeYhzYZ7/EeZkH8j3eMqjVUagdeFd
8qexrHCYDBffd8gGVnRY9FiHVJuQ5GxpKdelpaxPYKy51MlSTRNVElsafuUzSRUz
SbpICsklrqVQBR9MpA1BMKuRMbQDcsIBUGMUMBMoVIHZVNuXfWGdKDcwGM9dVbk5
KNGzpI0z6GTGuav2STgG2wP06AlcE6uIxFnEAEXMyJE4Pri2GjTMdhLrEwvDHvvM
VTojkXQfwlIlU5pwsJKFWYWQrgDRQSFLOkhb/cx/vyEKw9DjxwXiClZ+4U9kGRyo
qzjjPbjnNZj6odFIlOdEgqDZZDjmTjphmdW9z6axuJC4V6IKkxwsxRKHeZ+DoV23
gCNAH08l7l9f1fwDL+QExZLGE9Db7z0mcytnhKMrQs+Kez4WW6pcDFYcZZPcl/Zq
7Dvc7tuup5OsRIT88E83V7SDpbnz+uBjMQud/L8dpaP5j0lwdFZblLd1BWAplYQP
NGmH9B0J3R9zaNGJiJrv9wEOBJIMZed9YZbu6tD9ns6EUUG1dNPqiCpnf4aZd2me
7WjXMFKAn6JVVIoy9V7dE8kezXVcy4tFGop4GSIbqilZ1e4CiPtauNyqH6Op+QSn
t7zr8GUQ0aI0n4I/okTzpcjaVUkVjnrTYxY0aiTOETxlqKejiz0kFNdcGb+artV/
43LQN+VPC4FZOk3eyV9kbCVd10+C+m1/CUoeJji5Q8vMqGNM1lUuByo38HGRg+Up
T9V/dwcHYgpwPC4day3/62KGBSa7imrINgt5yIWIDy5jzxMhJN2ofgkLIdO/HT9/
KD6irmhi+GyriMBQWd8I3xlyxT1kL5eCZPP3hMcFEFvNURlCKkKMqlCJBFWTqsb7
PPwa5w69FVze4ijg2VH9wQiWulgNBIycdhTeQ3XvXMyIv9vZ2Vi2oaiRsUdha8OU
EtC3UcTOKu10Yhfr95SCym2HIxbrUg0eODkAoz+UyPtL8C9bd2yp355+BYotNUSN
h9JRsT2C3Zvjwb3HQbXKRgrz73nlW2hMqSVTLHMzkcb8ZQ+WTXEO0O3c73NFlKiB
FGbQAkvJIjoMUDaH07C7I5kK7zMKkM6rsGLRRqFEplP4Tcvy2FycZel13hODgJFY
bLQRYUFkeAMNk1DZrYJN3WskHW+KbFk6UxHGGva7GDzItWev6VBFDuWfU6t2KD4E
NglI9rwWHV1HU0gn7N9OjoLkxfdSJfvaEroRrvp8Hk2DKlxhMyPczCJmXu3t6iUp
1VhPjtu+sCMqG9jHlQEe82wf5KPc0BhwrzRkODJRMSQVMXYij/C2IAvIFoQaoQSW
+RR8KqORcYTVIzAaRzIgtlsuNiT9FprlZpcTxcKyFAXYCYDxXkWrfq7f2YcKJzbn
rDq9bXYy0Tuw5yhT8ylWFpj6TngN1JVQ5YtGbgwwlQusufFSoBd9DAEUnQRhlyKO
tKWM8T/gWXzFa6rCoYAVkRJQZYc1ATZsSQshKCPnXN6J5c9fJSu/JmxmU9IIUYCz
BBaaD0JpxCD4A1lWhD+F75RBCnSDDMzihyUpx7tSJAO5PMto80OmAO1tvbDRdhpq
HYeaiNOH7VSmJfBMBaEc9WiyP4XAcH/yvlB9+JidS0XBHXl4heAqvwnOu8HJrYgd
FlPToQmNkqpHAQR3V8j+HjMdyZ9csSGmmRWxIhetMXUa3Gmv+VdAWi3Stg81Zzu3
tjJ8OqpukZDhyfHlZzwRzWzteIurBNJd+kW1Iayj5/2JXFeodWJ2xSSZ3YrqsXX4
64qsQWzv6Zd+eHspHgg9SPa9omhDbQE9yvsxl45L2msHZ4I8hJnh7zTsFfFlFs9L
rIy7XvXlcakvE0DWpviGcoYa1T0uvlgyfi7TdzmyJEaUbOv7JDDiM6c4oZvUt2FD
sCvXGkjgBUDu9VEYfGzcUbAi+zvGvdJgYb4A3Vefgavvmg/X6n4YBql7c+VscC4j
bJXBYBKVA2AiaGn4RO964mA0lkjXX5TTH4zxmYjRF+xMP55bw+YOlgEV5Ig3gnpT
QQLSAmZPAjya8UbHMVYfkgn8xJ2HVk4/R61fBKcKTZzDg2QIEg7jfLX3bTWWEGMu
rDeQ1OBoYi25I8tFaLFR5eQnOV8N65YD1dyA3AUhUXkkUmsWvOApYENF0syVSnZw
kvfQmdRQRRNdhglRF5Qe+knS8px9AJHDMohZxYmmpacoolZShy2An1/OC7cSdH3X
yY+Fp1026uyeNfeQvPpzqYLYjXljEkvDv8c1Cg3xBkIOiQuSEVInwDoO2+e66G/r
wOib9AUtAvtPZKk08buyHLglR0/6t+n+w5bRcHJmpoZa+b6XtdOQ2a9LfwxdwvXq
JqehBacESuyG906WrDUNsYcs0vZ6kWQrKFBYvz8Pub/Cmv9vtIChTdJiwA3hKM4u
/pGtTYTiyMcuV3TJClHKmNz9c58B/fkzwbfV6vbarsgqwr0fmkYHsDcD0JHy6FtL
08RSprBK3kHC/KwX/NDv3oNIdsVaYhaz74tRA9hjVYZ1AHkabrAI2vG6p/D+aHPE
R/W/Ybj7fYfsdKkA4nRd5tkuZA2ptvtdPYju8YYqwjdc+xYeUaWHeLyqMuYWo2yv
DIAd9aEkrsn1JAD/Licnmd/pv/zaMksr6F6ZvlG0WX0YanfYgXtMldEpx+FFK0W1
1Iu5Wv4xb40F+TXo+MkoPwso/72yM2tnaVXaMai8PRHZSPqKmpty8WjUEJmq78Pw
+4cZdzaP/Qbnqaa+T+VbufOwvrnh3Hr/RrRaJjy1AogmANwGxbu0K+YwOS1GAwtf
SenwWcB8wbgjndEZ2CnhkDl+QXgHMwwJQbiS44n/GQoPNu/1jxQRksSGwCoGdp6E
rgSYCV4umqmbgE6YiKB727Vx3W1r4lH2/8IKXhp8l3mjFIMX2B47J8KGq/QZbSSp
ZuUI++c83vVwp0Drj1FcEgX7sxfeESMeYMem/Ha3ylUrKsi+M/EW2gvCsXJq6fyO
IEG4Y28jkGBUJL3f1gJ72kukCdHwbHc4foQ2cobBMvDpf5yRgRYNvBCWDxsF85Mj
4pjLO9JxdaKXAREps7uwpwVEhjIHGp2nzSMPTp6t8vtdpC9wnqvk+ZnA4Em7YZJ+
1wVabG/wEij+gOoG4WyYunpNqlFytxGzBF0va1+yYhG0aRiTY2737ksEfvtLH+68
xQsGnuVjrazc+eH8YlH/jpeC/mzQPWMz7inIqK6KQSf6ump/8Y4AgoXhoJMCyDy6
nJhjOgHWQprcGAWbW1pDMFnW4CxsbcdHcGH1JMGzTHvy5PFT/8MQIBZaJR5sYyaR
LTR26LVhDQpn7J/sYHwhXZV6c3FjZcHdMLFdXunBpDzkm76HTtSzKvkCft0yrV5Y
oTvUc7X5VMKEp1XfRp5ZOv6s26Uprk0QPmtZ0ZHcRpXySbcWx+pV+R83W1Zun/wO
Eqo/UyeCBwOeLQBNP0hSMoUOnxU4feDxIxiMyERqMUXpfQBH7lWIs0BbFyOSU8HW
AbKYCY43f3zi65f8SgXynOMWbUE7zix1hI14KCrGx6qLUTWNdysPg3QXFHNnCrfa
MqVdvQcP9jiD2jPtwO9VYuKfkYFAiZRXXUWNvTgErggd4UV0dLaog9SyMzU2ypkm
ZgZRZjtcAeaOtj2yk29yC8A3qTweemQnuzApr98DMn9Pq4S61epG5f65EE9n5Raq
KQySi1OQmJsp/2XHaDZTj3iururfCT8qmITq3oAPKlZgRnd0XDewDGKOwENe6gY2
T/3rrfbQyiphp+rZrjRI6iNwrrrMq0KDgTJg7qZuWVizZYCilHt96WSgv0Sen+aC
Pr5pcQxraOzdK65JEa8+JMD41MwkdG2Im4XrIURbJDghldkhc+V1ZHrCS5zDaDUK
+HEHd6mY6Dg2vLcOnDmaBLJeiFdIwmTFLGmTQS9yfuYLCn/NgXKFkWkeDAv9YpHF
S8FzdNcUk5TTApNoYGDrKTd/5YXWrcSm1lJnqAuE6j+vfN5ISkGuOrkP9+yvb91b
vqTSmmmKro7C0JfgKZ4kSBfFPmsJcAIVlfckiQoxhWWKUovsXm/Q0iXmXEGiCn7+
stFNEa3g6ifrSJhUZjlOQ8TtKgauC8BOiXgIQBplsksqcXSDvF9slG6/BFVi7J9U
v7VW/PydpN/RDmJlhm+T2MFRzs3xy206iPlMZ5152g+HOhcwAw49CwmFmwT90F1A
b8T1ZfS0Dq+eVXDoTZLWCISfbCoRD6K9vNxmPXVIVgTYQtRkfyOVNHu4EPij3Zxo
cqr7bPirGtaTA2TD6aYnb3+JLyapBEZQpN8q27kvtUM6I8BTa23vU2G15IJJ8ht4
xegl5zfGH5zKZlNkJzWi/7Lzcr6BQV7IoskSJZiHaRSaH9Zabx9a7/rOFavfpxjj
YebaE6noaZ+28Rqp3Mg+HVS2ajXPy8/3+oJIY+fP1b8drXwVijNVNtgOHqx1rZDs
oqJKmIO+jSNAp6YTSO4Jr51ATRf7s1hF1lWo1wQwW3gw4ut0jl7jq/eSNBbeXbgO
C59WWXQGkkOjrVOgMQkK7iScycDO5Ra/aPylS4DX1DT4g2tRkyZmldfRLIZd2fZr
0IlOqfeuAKtp9YvbS87j4UcWPsItHIMbfi76H+WFyUXNRFue1zuVlntF0rdarSuI
CuOhrfrZ81ctx7mZcySJK9k595wyAWeujVvyfUyQ8dxmKvKbFkclAi2udFeGBk6r
NIJ8hxPWr/TpCV5LTWQL5L6zkEq/Nl7993ShlkNfuJY4Tuz+lyP1jHMWIlb5RGyS
YVCs81JuxSLSK4nUcYgWVC66NJ7t9rm5gocHMaw2ayIaQeZwxjl0aXzCVZmB5gJV
hGodWWyYn3yvt1AjvszHwOWP/XqUajXIeNjlehiUMIHbFS4MNqFFzHKDYcgLoV9C
PveKUumZizpi0lRTllTCxzVPBvjk9RQ8ynPippca2xwYJUABCsTUmdO/RwAljo8X
FfI0vFLlwAcwy5m241YKDOaTo1heSwgvnQwEm2RZjT1afW+RoE9K+Gwh9W2r0nd0
0hvEkGe7dFcAWSIK8bvqNNDFvkHyz0qfQwSTI7+KpGVnt7KkiiHbyt0RvHWk37n/
FhZHhXsGBvwYOImx8Ngis5U6i+y+iuXefTgQTB6bML/c4glTrVEFn4pkw2dQJwrX
VXgKcaT70VQgwJ9APx5i6UeZKngAWWrK/34l67Tj577vFO7eRSIdGvrwaTmeSg2i
sEXRSIecPOK36pb964VFWfKIg9R/wMopNQOsJVlsx08Fjk/BGRqar8KUHZe901Kk
gpy3uDDjHiAJMeeeTbuy46yTK34e4C4GOhyG9oMYtfd0FCILy317qnbALyjZh1Se
qJNn2N/N6shpXH4cVbIRhGQ4/DqhqzWXJ/X/oT5BixF3I1ckTJMg5uHWQUyxrh2Z
sbqwvoLcPrVPXHZyRoK7hrvIgEulybF5pmm5eGjAnwRGcwCjNiYCwDD28agYD15Y
9DOhUuTvTJ3r/TNSp2VVPw7N0VydHVCJj8FBS7N+T+4JP1nvGbwoUt01nQBVYtQw
+VrqeePNwyaSqA+fzXwgFztqZjgXR6uRU8KnRYzT6TniE7Dqke/3tuaKFbg2jB+X
yybDrSX1I6GWRmVZfgNaA67kWtj9TKNh2RM4Ev3SkDt5kD1ZV2n3FCnjwaFI5Adw
E2C/EWv91jGTBSo+ct2y2MbRpcUPuJCs3FYuZC2JH2Acjtz/+i8N5abX51hxd44V
RNWYSsWZ/ndySILfg+M7n4VhEwtmXvVh4JRbmgZc1e3/Y/wioaaFQOAucBKhERqI
3DniEaEyHhJlqS6DQW49tDb6d1kTnubQ/cTc7lAX2dEwIfywNQyxO78tUYhU0p9K
Vdy3T8DqTSQHfA3d82MYrS6DCGsKnzGrbCPmKO4RsANuRWVSEDAhIlC2AAdAWFfZ
Gx3G+IHZ6Z17pN6JbBnjnugZV/dmAF5+2sbwqXX5WUW/6YoYLDQNHYkf8T3fuK3V
nSKIZYHi15/nSo9uD8jdfK2O+aJ8b1vgEpSsq+JEVPph2kz8Wu4r+ARxC9Cdx2z6
3K/FglTVBC/jpitHZ9weFpr72QKI6vTeaEeBVLQcEWVVtp4NyrxV2fyJ8zuz0omT
K4zT6GM7KWX504lTbUso+1FE50LI7z874Lnl7Sxx3ketpcM84d17DR8rLTTbsdcM
1TEQ+wmog6KxOmFnWXBu/D8OZVGVP7ZcOTDStahKuTHxoOxulTbkWWu599VbQMA8
Zd/YATOqaBjqTp0zjQSasYgeLSn7D/5PhQUPVTdB7n1e/g3FmaXwSw8KyUSSMvkp
ZVArZoVaHdVm7qymTKQrHSJPwrWaagY7w2/NcO02B/0yZUwFd941AgnmOv6HfNWu
Evp5UiQuiQ5o6ZQokW2Jt6fd+53xDky21KNOvgk/eecd6MuBQbHDsHVwiu3+zQBU
mJZuFt+WomBXjz1KXCRgoQBkisZa1cYlhiI67QH8eGKS/b3WrY2EYJsoRs0m/SjC
RE6yiLgaMZzmBPOGIkcupBBzeaw03mcBb7oj/WwEuAtbdD2Nd7b8tQvh/+tv6F6p
O90nInpkfDB/8l1lA5kYLuHL3/15kMbr93EQZ7pv8JD391WzYww0XWbi0nloH97s
I5WNr7nAk18Rj6v94bR218PpAufrof8BRO5Phgmd0lJh1RMAMCcW1ZMxnx7m8EZk
rL2pNxL8PQiTj9DDhsDUL49PpUYsTwhbDHsXQRGgTdvY+RPtyib9wb7wcdMWdRel
tAmSnMGzK5/4eaI66NNbQ9lq7JTJn+p9cjqTMRqT4gZUb6jbB1BH9qvQEW4ipnyt
F+/KewBjL5FeCfPJv1DAzDhJMaOAAv995E09tbVNeUH30W1DQ6mbscf1/ieLFP6Q
QYs2H/vGktVbvBzm5vHKDop4pTcUFIUjKEJEhf78ODFfUtQUrk2A3MUf1hEfg/TQ
MWNOCffu2vlFZROeUHvSo+uLCLtr+4T6hCCZtHfMD31PycdjI5zVZqiCfao344N6
/SwT5jYCdgB3sk2BoDWWRDh+HBidMhgHd1wE5K32r2WGmX7BLOaNPYId9OSNQUaP
Y/z1lBjM27uIS3V17rmnmQrZIBlTplHqO5T15Qc8sHbVyyIRF2FwbZqsKFBWkWDP
dcz/cIX4Vmf+wTwnhsN9CL9k4+9+58Ke4gl9GOBf+6oJY8OfTSjjCBttpjdIk3xJ
63e+am59dS+Sye21BAMEDH0YbmQczUBlTbN0kfYT+OmijBI3+LftHN/DcpuliVHF
Z6qE55LkuNvpCHLc23tR/BDu1AXa/pG+jUn9GwNxNFz5t5/BLR/4dQBooASAm9vo
ERtxJNKbvfl52nGzrIMPOYEZKj/k66Dlj7S44wALz+xgyZ5Lv14dEvxOhxvM1mtL
E0hflQbfyotIA1Q2LnT6zPh62TD5pO14xuGPX7UYICRoj2uXdzc0SGRCj+oGv9V+
Voiu5pzAcjv3U420K2uZeGCEB0Q8X8NJKgqVRSoKpdGoz50lsEJJWgtyAe98pqnk
h6ZCPM4YZlek6zY3V0ceW7xTpZdrkjaZsNKNc4aDrEb6y78C1/5sOyD7KsEC4/nR
wrfkMJoI+of1pqjjguEOm83wf3hmVBLOUBGfpSmHyYlarI74lLHYOswMlYRWq8L7
UmycYihQq2mkIi+rI6jlqtJmix6zgHMSgO8WiitxAxfMWh2bdoXR87187XkqLFHo
FxvPTxnV23ZrnJRx8aHws7C4DS8A/4bZM35aBf3Yzw481Zwt/2DR+WIN9/2u7i2a
N1hhxFd6vXYnQvGiJYjafMFEvjHy70IQmobGTPq2qVZBPYLijUrjkSdzllrN4KtE
98DX3+/wXCNOwb9KeJB7P+8eD1CPR02Gk0aupVTjiMK8GOSa3WmM2eURWQE5pnzs
/d92BK9pEq63LhxbQxE9EbEBSUf7Q8SN6VWm5SgIm7DtfH6I3JBomEs54/FGtDp0
peFyP52vFwQenW6pmrXVTzXXAZcqnwxp9Aab+dg7wNChR/TJW4Qy+wckJFT+hWOA
8ZP8M2+35dwi3XOwxTq/hXInPcff0CJFPwPQVJVifSe887PJIs+AOqsSCoV69IeU
p2Cq95Z8LvDJB7iAu/usw1CSNf3qctUPlJMx15GOMTVwuPH7xD8iFFL+OCGZ6NVB
2xYnR+0lZx5hT0BO68OYpz/7JIny5TNHxP9yJ1n5VmdBLQJhNSUx+jaywwHqO1mC
W1mv3ZyvpYV0SEMq6dvt06nA2nNunpmFyCt7kYmVYe4xYEvvEiLLLQ/kEFvHeg+E
r+0OrVz9rTewG+WMyMnL7pgb+bxgN1yCZmprdLnOUXKwYg1rodSXLKd4Zd1q9AV7
e0ieafXDh9BPl2c4AZmLZW6SekLvo2kweNWtS9Gknvq9J8lCCT06E1OFuvwMG7G4
dJ1HHHnnisMDbZqZLxSLXDIZ0WGe09LDd5juoIPuCW4OdpLbS6ieIFqxEyihnc/O
WpiFDGVR3r2GVbvyZFGk2acza7O4XJ+TDqJrz3C5nXQbs/lz1uYcYdydXDT7m7G/
vSsWAYDDFhzrxAn9jNDqD54F9qERGrkDRXN/BxglQsSVjH3/HQfjXJvmiKIFmsWG
gfS9W3/KQZdoYu89LHSVea3LJoaGc9/EnmIOpYvFXDAEpqMvWeqCMzZmKwX0R9WC
L0rG4ZZ8vlPXamv1KqSmDIKJM7+RuPVm7qeRtNDCRGevfnO0QGoBSRkpZ3rtLY6k
228kpBD6pGNE2KwV5ykDva7n9A1YocUMAqYXnE25nL4F7BBr55ViPGxI+zyddGc/
R+iFAAYODdL+JQjFlmePpZV51ttCCuUTZbC4hEJ0BIYISTBcjqnVE5dy0GZ0JkE8
545wDmZqSuBV81WQf+Ka7pnQ9XFgCnIW2lzkMoV9QRqb0xEccj3L1P+CQx1jM4TU
o3qUA98oLH5UfOXYGOHTjr0aghgTEBs4Qapf2a8XI6kBvA1qENqi7s9eW/OYo6xB
CozWO6XICodl5tlLOA/rkPjVpWivdJMDunwaSx0ujYV/RGhkkPSJCNq7fV6IevSe
INtwgc/c5IrX/06SM8wosFd5XzkfLm/ebbxBhhRqVT0V5YbJkhZx8oEuW3p1fTtj
LvapXVn9vEs5fhrpxERKYyqWKtamaMA+Z7uthh3JREeNNbZxqCbaD19GRT64Fwe5
RiubHRSvBC+1iVM9Uoc/FoHM46lU2NeQdMfGp3SG9Tb69HmO2pcy705BeCHdllBr
U+kmlFYq3AqQ6qWIlh8MZmP0kzHDUpVVuPDXt1YxCyPeP1Cf4as4wuNbXtPoPc2q
8PGjb5uqG3gtVD1GBB7Qb+iWJa1uw15o9Lf6SvcruADtVzmZPPA5Ofpw78s7qxLc
hUttkioi8+V/OmEXntM1sE3mcUuwue67IaoVeIiI3qtBJIZp1KR7QiXhVv4bMolA
zroiIAJcfkU5dpYAj8bIp0fap5NT+Bp6XLHAktnJOa/Z5NWF5XwSIrhI3U0z4vyp
DQxKzp8Mpb+wlJWtFa/jkS+hhplqGdnSRg/NMF3XC6SB2DfZBEOpFCFkouUwNT/D
IP3WzCHAcgJ/NQ9fgaAULS91VDsWtjSyCYpXV3d6cbGqdByR/ruTXNfJFInzqi/0
qfUkyU3bZMsX7kba/LHC+kLHKhoLMbLicQJRYx+qLQRi/CLtKrHpQUxxaMpMXr2Q
8e1f8udqWDeDGAqljRRuCWHovzI/i5rxZoUi2BfdPds3toXPDziRDKLZ3nKZKIe5
9j1u67Z6pMbNz0i97+qNUeWJ87K64qbIgdBhJoKMFdzQA9WIJTHoaJkf11Nl9l+g
aT2af6PszTE1MBjr6bPTSqFtGDVgyyo2YtYaWfacdoIucQqzsGaI/6LpOS46h2hk
+KJvNY9el1X/0WiH5wuLmxrxSWqRjxhUr4W2Ff0CZ0+bk1S4tqS065Nr+455N5Ry
L9ZQjlfORwmosTEd/6uR0X9APq1e8RkcfxYdihVl1jcahccO2ZZbYMiNZ8sH3ifN
6CUQ7hWwb+Qp2fPIihgMdnnUOwlFqRaw4/tEwHk/uzB8PHzUSge7QfWcur7rNCgp
QTU6G8wZNNb7BZhs3btHnt69bJZlArdjPqI+A9gfXduvnSiFl26fDUY1H75wWT2J
bY1a3iQg/+zyZA9Jyu6fdp8Nn1tZgWuKy5oGfcu0GBNUrh06+dVt0VSjB0WcamRZ
8hyCW7/puYrJ3x//+YkdZHit8QFfdUd6Fn/z4Hte7ozVh7gtRT7Pggw9lnRjPOp6
xZgK1Fcv1jVPCjq4QP8UiG/7G+ob+uOOhdXyrrNplMPDqZklkrnosq/+XwbI4SfN
+42Z1FSz2bqXSR1RZWw/pyCAR3Usg+RBrzeIe+Fy9CK+iJ0zjMglnnFcg+6fNATt
pmbvfp5coS9F+iszV5ezAHiLeMsa1nBdGRds/rI7Rb4sEjUAeUxi8orTUxnMCldA
oNTwnMHTUNesjQ9FqAf8+A7kgHTIKa1Sxew470b55kbOYUiY1kO3um96BGmhTGOP
Oh3rnMq9POYs0sNj6I5m7HTboo//v+C4F5RADBP9/AWVd+NTusbsZuFXnRfQ1e44
oflj4G+qXMvCaqRTvWm7NnZrqRWb/G5gEExZOajsjRmmMmHQENuf0yBEfvzLAnZ2
yqBNwmYZaJUnFTq/V91Za9vUyfAllCcPBCArKgjwf36G09AbxDW6brgdsGRMVQs2
5wYN9hc/tzImC4aAVKTtFGE4Ki9Au7/K+scO17BxTH2Y6om2hHGYCCmac1Pqe/a7
PXQx9yhNh3eEV8rxembXKvzAQ8bl/k75rsddNeK/b1mqOiRQAJpcmKZqxq9IZdNv
DGrTkBPPzXZtFmwUM5GUw0pnJdITqNLm0iTvUEJTuSS4jgvFE6xIMa6/lRdDpm87
VDtubT+eY9BDPp7mP88Pnbg1E6lhybpNMGGIPgiJr2d10Ocij6LF7S/L/GGadpei
3IBL79UEf23iRj5ODOf092fpvMUfmyHiGrrvvD953qT3jQG9IDRKfblkZ8fOUTRS
YMsUOJ8O6No2HnCneNykm+Rjvt/v1KdG9Q+hyFIqrEdLvo8uxa3iSxmcQ2IgMR71
NqYpduqcWMp6GpzACYluPLe1CAb7DP+SAZTGvIyHXWgpJ1gLglN5k8TSF4sJEYXI
7tmgE2gSEc3ynY2TFbiRuOhAkUxIOtpz1agdjvhSo91QolueEwlmTbOx0G/evwe7
kbAMa+yRjACMikpaAiLAZg535DOTPUD4ou/yEt4+Ge0347zUZZxB+eDL620dI4dZ
p2NdxN0wBhrOCr9gqgbHDA1+hDvky7N7aiDDNAlZYsfRukvyHaG7U14KnIMAQW2G
vUjEn//r0tGkSCcjp23ogwKltvoVnGas+9QutbhE/uTYH1STCbIa4sMZKzVNHpYX
VEUEc117GxziE5gn20ObTS4RbHycwTb3qjH02qruoUA+ASp6pIdWnNSrL/LPjUiY
q/Av1eRBM6Dwg2UMRNc0Ya+Qc17MxMIZ3hMxEQMJRfkBk3p51d4h6kEMx3QduLru
6DKUtEYKiJA4ItIrCsdaTGAXLwEaFm0aBkVvPpNH6IVybKH9ZsuYDSaF68g6ipvc
h1DCnURL378Pa+CLDBKozVXK5BZ18s9uKNFry/uKdeJAFCLKmuvTb1IdmF3WU1c6
zxA/W18vhXfickwBnnGyg98AXW5UlzibeM7dD3jVb58/yTtQ3019gEr/3QjZhRzJ
NMZA9zFu4vaffYgyJ0neOqcLrpHwaFp3nGCmHDS1L02Q7J/YbGMwPcVhdAow1wko
rz6h074g+pTZkQ4H9uIbp+dsDlEJKKsgE7s+nmqzHaOdYTLt7FpXQ6V0J7+UGfbs
h7gbyovVfnncpxh46gAMHJ+o6srvSXSZCgAVe+LoihmD135krAoObhdqe2KMCL1o
j8SJ92J4yAhKxnjjUZMzrwnEhEZIdHsOL6O0RrDYI9tRGDqDA/Hiv07EfEmX09cz
o2PsP5BtceXPKt7l1hXAxqwb+GXz+5j9wbgK8QrW3iBSwaqjvUIw51ghDn+AbNjG
6LTnlrNRQjfi3KzyF0WEoUX3FfzXIHJa6Zdn1liU+wXkpM9BVKwWJO+sh9lkPaPu
9AP2aNPpHtT+srQmwmj6aOFUbYRWSbAw1vZ1K9WTXgtlEs3pRqf9rBXw0VLy3mwY
vDQSkyUPuGabMinnue0Yyn4dcmzMcmvQsHbvwmgMMwg4ET9yZz7lbvwk2VNX4rRf
27J/+v+DgHRuNJFpwpZKEPeYjMxlKRqHeI417EIwJfssw3/j9HWF7wZV2sDosTdv
R/ux61ShlZ+XPcyjXrz2HvEShFh/8VZ3ebzqxfp//jxnw9bE32znEPjrwa2jj50J
rehTXpussD6JtNZlp7U/AiqiLgAbiP//00WvQbYCu1y9N+140r6PDogbSHG9Bj4Z
zoE6J1CjUBDHO4R+YvRKHbRyM5+oUi6lfdJr109qE3bkibvVy/2+uoL8f+50QNAy
1+0ZNzBCMLy3rIUz5n02Rw3MHu6rZUHHtR9x3BoZLcDkb0Fm7v5O8A4vvnFV41Mg
aOvyaV1yBIgeS/wOXwYvF/aEZRhXqks9Fm/No0EBHGe5x8OQRvJIbuy1oY2Jd+TY
n13Zd8EB9NfO8odvaDttyAAsfJnp5jtWOfNrVa2Ko/6eVD2FHn0nsgYSzf60/U3H
SIrdYbx8jBb/SsuJRpDglpjDvj8gEjrdO48A8n28b0/UkL93FzvhgJWpPIa+yab9
TmyAai8uZ1a6SzhCI6sWp9ddS6ZKtz0YGIfkmquaUcL2ipymjYwQaOsqtfgi0z0s
/fdGm7gTOrEIwYg87cF2pGZwOu/fVNyIUEvWB3epNPdIuRHSkGGRyMcuXQLuAjoh
lqkxqp6FnNYqP3PpXKkipenttMeYDv5W6/FKWG4QLsj1wyI/TIJBM3eNYxFPEUQH
BqU4CL3rVVps37wDkGNor3C5MlInPBq3lDQUhhFJl0w/8RUeIVgG0pj+TvILAxsz
+CAK3wscY6UgeHzzVNwvykEEYa7A2dugIAiYEpGwODJrIyCSTpI1hlfROGjGiSNV
OJLGwqXHCO6vSGhkEuChXCZmILGYU6YZK0KSUTGhea/fv3XH5I2JyNY5qSCG4FH1
sryPuFRL1RSo+KTT7XPVbol/XjfYOaA56kejAiF4ByVBTAn0iJId7IqE7yfq0l0U
vkcQfpkJNs+lpGpGwVC4MeBi5CJbx6SynfXGxZ1chge5TGjeVfz/OSSJxH5lYXY/
QXJL7IMqm1oY04WQ4nk/MEbgo/Rkw46dOx1ISn1IjKIqn+xIpWyyiNFTM0MGs2zF
LKa6yjxyw1nBjq82jHbAvWvDGyWZsA8Slk/VAB8VDITXv5i5RYh1x7URi3NwEFqV
a99mbC1u3GxQpL+TDxnn28YWArqvswCFbveomn+bB2RM7fmkoAnaXL9O1yn+/qlS
v9Ah3+jzSYd/DWyYsDmRY7uUdrNvQ3LqsnB8mOsxYLmwdPCrwaSkfq21Poi0BhqP
jNXSaG2Ugsm3pPA5xfpHKahu/8mLTQjEVj4ZjNtLg/NZaeVTYxatFxBfUgmJhkGv
yodPlgn13abMAka3ZO628Yv/VxahshwxRJD3OQ9EQ0X174yd9fJk1BhyBO21nynY
zSO1zlBi+2uP9CIje+Gdf0+lB9qhi9toOxbc1aSIYnU6xl25SxgsQT3Z7NHbz2aX
wCE0tyxDVa0RSPbLJSHyGSRHjax0adTuDBvEhD50zZay6MrzPJrw5+d5UDdQmF/A
2OTVbpVC/DQq6zSEM42wcu12lNOKkKjWlFobzOwRvbnQcbg8Xu2ratHZdaycH0B+
RJxBPFg4ec/twIXQcYYTuwx2O4+3RzSb+fNlezoY8NMRPUvFfMqftN5g6whHVHho
R2vSwhOluvbs46IkHlIgWuReCLmvN47X3wJpf/XufLpF445nL6Z8+aZRhNYGsyq1
1igXq6UFe+WJRH8VP+q1OqgjZXNw5MsY1zZccdBjnboJ6wwzEfKxrm6JYNnL0Pym
uCPYSVWM0gXorBd8mcXTq0S4hTrRvMPruSexKEzfIJ38N7CNqnjozre6u4vHG9FW
iZG38O8q/XunvL8AYcqLa1AbbWizcwOdMo4z9t77nHzpQCGZENUjw27dCt3oNOFG
GwH6doBu0/A5jqdmQ9MKh02+m+UmWzxt6iYyQsf3TvqWtgAa9YOei0lpjt5Sz4DW
Ssiw7C0ERyLtiL2RYqFKv6qAKZ92Mf+DJHBPKPW3uOFgWtws5XYXKCAOC4qOPGPi
jd/efvanuUW+aU2wv5XQ1AUigI8Fhxr6UbjIywVWVbvoB6KGD/Hk//ZFQwQMrGX1
tYfkrboOlgq7ggCwPRJiUwjud+5Wf8k7DnDl1Myj8Vlq0G6wTAwPXn4+epyADmcO
/sCkb8Ln1gs0sruJ0Wq7M6Uax7DVzg7BIJgXYCgNEmz0FBEwhgKdTXNr1AEwLfjL
lpL/5KoA1zg6Ss1IDgUSgT+PVvSdnqOnyJuAM8EGtelB+QOOtNDvAedUN8t/frVR
VLWR2KJ+8NxCP/dfuO4VSXU0UJ81VqplRxAPHw0SqS45+oUqvcnQ9NMczRs+cAVB
REoYsKhX89fFQVny+P2BjntrE6lkGggAVB1x4l9gXOc57ldR0Bc+ewh4fNNVQSHf
5ab6rOAuJ7Kl1FOQxSlAXy6aYoWPMV7/ug6jFuQSJlc5OiyrUx1k1ZhwOUwWJAAA
YAw9vvJwxf62XBgQLVXwzVKR3f9mJMIDO+8dy+N+M0xMenBt+uA6edTzruW3/o+W
98C1dpQYF2W6gjR8Df0I/Yey0Rt1amOF6JwnoKaB4Oi69HArYHGC4hi0cUiYi5z0
F4KeYWryD8PIiXt2Y6MDOCAK4x9HSwPr2ZLmZKQh7ab4xtqaR9GJmnvBCmBb93Ld
02zNUU8pWAMA1C0QsAciwUTGu84e28xjfYly+7Ht2CJKVerXIGl05C2BQNSboXDU
tP/UrHMZpFeYH9D1/kAS4Rzmx76SFmHfSg5uYXhvm8Jr6i5SG3Xkk29zU++ySrRS
Y+37ebamd6vNK39OSr78zmD/0yuyk/SIUmFCMv8f96XNhhw2ow5H3fdKIHezAVbV
H5vsVfwbMWQfXmVzZNXNZrOR2W9e/ZL8J5VfX69pCBW0iw1twDrtTBrYr1ojG63Q
sHTwiw4F8ZCHHT4nURvRPNvNI17UjjQR6jHrj46wcX+QovlvgqDi75QWbOd2uJCe
PLR0OhhaloXSUecIT+6/dZH3bqxt1XsxXyG3glRnlQDwO9gSJ1q8HesKbgCQHVUD
KwLJWTgSbG6S8IH6Mt8QYLMnBIGDFfpmCfXlsebYzsV2r6vDBuU0pz1kME69qQ8d
GnxGU5Sr9sIvdPJACMxD7Oi8u+sY6ry099bW6F8Nt78whm9MHeXBMZJVO28a4Hxt
BXWMwEtmKvsb/Rv8o237OeXolDKZz3NTYDRXPDUkaZFPdE5W3XYTJBdpFtlfVEl/
e+KhVcnlTRm+tyoPWOAjgNcf6HHSq9B60LXWY3N97mNctjHouH1tWcEcQE/aXzf7
CQXMCtnT1IfD1K9lsFe1gFiU/0PAtaRQINn8pJ6PI3bwrdKY2ovSSrVZVIk3Jr5A
T5ax06XPO212wq5H8Tb936yXBLQLulrt2PUMF6nVeveCIKcTVbB/cX2jrewHZB9T
vVQZGtGT+WlQrnKUhZjwVaoF0Vvf0Wfb1U5cQ3Y/L/fq+MgkhvGaiU1oTQszNZn5
tncAF8L0/xsIaCAWcZcW8/IeAZPACbNodjRGHiGL4D2ScI/3fwdLRqGFaMT3D4Ou
I8lFG/MDeamiqCA5uRFPUlcoiZvvyZCN9EqNx0bP+gPXliqYvwcNdLqF6XF6xp5I
m8zFxcx8HQ+fTra585Qq1Qw2A3cmTppII3nJ+d8CYYCLNSPHqsozzStzdS+dcfZs
IN4+neLsNkcBRNwe+rdNX4m2c4+YXBoyu9EARiYikQH8KRFvMuUbOD1o61ZC9NcI
01pFT1wJd4U5WQSkaPLP7M/zg549PyGIhLEkVGTp2lGKO2u09EDRnItzFjc9jfM2
Y76LWcwOpGYcXxOqfT+XsGBm0SUx1ow14lnt1rUEgPonurlYJbC/paK3ffmx9kIN
I+slZdctwAdff1RIEw/dvssuHOaCx5sWmeeV5EqTPzTvME+PrsjijH0zJo9GRhKq
Mw4j02jfHOigINVBoA3HX6ZYNFjp3ZehT/tB6jv+R4dJ/ymJxXJxpVnRLIlIdTts
7UY3KcUoCV5YM/qw1Zk7pRAa/js7IrL4U0MDbE1xrntvduDX5+zbgBQHU58YNxGv
aY3YZaPMtuZQK3kM/RoHrnKxHGAprn11M9qfUOL6YJm0qTWkHXfuvZVl7zg9Y8yv
KKIdh83uNxQp5CP4hKygYwZqhS6S16D37khlrvV866DeBIogTgnU5UP90HrpDioX
Dpxkrlf2uG1WyG1xN6Nlh4ZFGU+GXGPLH87TmMi78q1NWyy4MPjcDWlqs0sf4lng
USrXlv9lQvjf+iXjjYf422zyiLCwCXbP0uSxfMsYCnAmBnd8QW7C5hDrn/OVKVgi
MV7eAuE59o33IMXNkyglepORORC11249bqsx5e5Nw8eOqCaFpik3C+GTpPTzMSCV
nuohhshfZi2+7wb3xUatyyBhrOWCiQrmyOmgYMb+gPQO5rgx/inhWp+hLyy81Nkt
w3nxlHRGSnMa/Puoq6P3jVxdSLdfeQ5wg+MKONjHOl6QOgI+ZRok1ZSKTqmOPtaV
AT2I076DVCV++s4nmy5e6uTZoT+bJ5TaXlZfTiEb7fiEmIeTjfApU+vXwz+Uu2TJ
gjEOfP9jrDiH1CQT8Az2lbCWcIfE0kdWfWyshAFxdIze8bNeYPa6p35PnwqUgZk5
RIXltec8bRBf0bIo0KJ6/Y1CcPScsh/h8YzQds7HawwP3ma+wPEpIehTQ5IbQaMj
b1PaD93rWskSvU6RKK+XuPgeV0xeiMQyDnWsaLOJhaU9ThUVeLtcWLZeLT/teRCV
elM7i7sOgEViFRrDGoq5e8IkLdjOTefJBzXJ61HUOoKpZADeH74TIsqk0tg6Zvq4
pueItIBOKcGw7V8MCQCtAZJB4lSxN6tCcVJFl2/79P6iV2gg0v05hNeVlD4+XuoL
lKUmVo+m/JDmRrHXJJKlRBGWQ5R/7JkCTgU9wF3edX53S1yZlJrhytwCwDsr23NZ
ftjzcfD3EY9ZNgBcMpQaRAGOCDSawjvWB3lw0Um20oF6X4VqDuAv9yeYuZZp0zWm
ClOOL3LDYZFR/DR2qu6GCvVBNB2/jgDzGp62CygWDR3FLGwHv/m5QXGfRHcGp4vK
HUIrrNhdjHFAyeB3E9wCkh8LOO2A7Msv+XVx2ErhUpTka7zIqcQ9KA6pw7U0SCoz
1G1Vj1lsJb6OmPAYUz7X9Z42Vhhe/GUEMCTm5BCHEkiUoZgRQNrm0JQ/0HeavvpD
CmeakNTAHdBkcCxfRXk8t6ENVMvJ5rsrWXvsRPgatPdC6zW30Ebsn1rD5l3QDIXE
BERNZ4w1d7pdyhmQ9nroUY18lhVQkMeCQT5t+ey8bWcPEg+oM6XnJMQdXAeHEvVv
VfXmTD6N2w4tZvjtl5yHrp0DyEPbGl4I3Pr3eIWJ/NSB89EL6bdIhplSuow+Rrlg
fD7/OtCDeQc/xTPYsreNYr/dhGgNXHwuCKUsgMXYRlRv+RuhCGQHcMt5LtnAQBT/
pIUDlpdZPae2i7VTwtLza7IkNLMvw2Rnn/e9d3LpGsBINeO2AH0YATX1M5iJHdp8
KHY0M3JSSQwgtA3kvEpP2qz1Tq0Tu9m1T3Lycah9xr0YHBaa+BT8jGjv1V/dIZCA
z47ZfKNWBpmz1pqkEDfISwgBeeclUaKqBO8+BCADqj8xW9Yx0GG1xXQU7CoSGuif
bxEBRDwrZT7zTLX873V/K6x79OWWoSnuRHPW7XagDAecL7WgoyEEHwZM7DeSHmt/
QYktXR/DZnJkpgoYxCsJP28okpzApjw8vzmKWQ03MsecsAtLczWhqwu9i5PReFg/
mAS9nGVjUVNKzj4RyC6J/BGLyX+Qkd7ESEbdXEZIh8Uf6UByBwC/AOT+CJ/3kyuU
FDdL9e4oJqTJdQeo7V2RT4tqKm6PCJ0CXYrOn+R+6yylL3RfyGhpvDiUIh38W6KD
kxPRfxoAMTpfyQQIr7g2rOlehcE8MPIZsq/ZTxLGguXsghQeGmHSIuCzG6lmGLZ1
p7biogFNpfJHQ0FrUDZ7ZgmnMWO6LNeIRUHpJqrO0TVb9VjjmtXGL6LuG4RL2H2X
l5L5adMhS2KNHUO7ir8sEFknmyCwjjLgRHmjkoYbyC+VYV4BEduhKfMmcvf+x8AQ
zAGjFNm/eKiFLkATsZF9Z6n5KsJDiWOKmkBg9rp4RTJf9n1FTVimIi10JduMp0Sv
s5xtgV+YtSE0JsgdnUS/eMqBtPXPUrLbf+eZdhPHUAbOZsOlyOLTqwiWCyAnEVeh
lTZVE+aqDYRHuo32Dt3GRBtvznksoINAIEmV2X1ULaMJ0s9h6WaWqj0H5Y2W0n+X
4vchz97eFkNL5hmSr6ixKeu1BNMcKAmO/F38kBR6+P7LpQomjBDfLZRRKKUUl4ap
gGlJ001zM6dcpCJaBLr+MhXOcoK/41f7PFXcDh2IAG1IAXmaz9KZotz7LLUtcH03
aO87kL0XafplLeUCPwStk8EN/L2L4Hy2FOyj5eXNkA/DWzKmqGHK0h+KyBN1ZwaQ
yGJJFDVm/uUM2iSvFjAOK6TjXfA8FIXHQv7F72vvxNjxM175NFTMNlm7b8Kq407K
iaa+RA/GL8cxFiMUe97mTFjoTSAGBTaLEyOgmodwRalTRsQ1f/bI3D8Ef6nrgJUb
Q4/n81mYDAqLm2RdvJPZjV4knCD6T/O3yq9LUeUnW43uneZCHXRt5ZG2THGWJJaR
EQJC2Z5riq2/P4QLkUCmGroTmCzzii0YLpySTTM09Q7ZbYIE976UnqlHol7WcIpD
NaYfLuuckIA87mfP4pVF6p2PPtNAgnk3xmyT3TKXpFs3EH85UDGtSWsfPU3s5+vv
vyKD7vtb5/82MiStNju3UELUQqhu0Ukpd6CWnbSJucSPvjy5aHej/uHbFnOCRIcg
0lazGQkbtQDIEG2cu+ClRmsWT7DM26ULLoHmIwF7C6MZFVNU11+hdYMroR5F6m5z
7H4motl2a2lSwh7EnDDEV+ag/u+nsF9dgt0tReBXATPL7YNAQZZCHFTFOuDwoOwb
2QykvAj26a7uOhpeomr+s1lmIhPGF37MTsDzsYviK7VYquCd8oY0W0sXCWVIcvfb
TKOlNfJ2S/laQQ775U559KMXwj8N9C6WvVmzY6UPFr3WaLgBZTqta1Tkon6nO9xc
swiZb7kRtHMwg2OxoZ1V85Wk2tOBg2HDe87rl+PaHiwm4ai/8gQUUhp3WwAQFllr
KZUhyzOuKcSn568vP3uBGOnzaZ04Xm6i3h4yOu/pSK3ERNpJEZn8PLcBOZ2urTQx
jhna648FQRyEL/yQWYylb4IY43+mbuIFpzvH5efYl9LfgydKoIkKE7qNf7X0vmMe
j4PuXrpSO/pneFBPSzVfahhBUYikBlPJXt5osLmb/PsY0zPRz0uc9p+jMIB1br+g
tz/FIf2RFqauOqVEL0Lr1YdusgVq4K6nFYojWMPKkRpoG+kzia3SxaoEplEEe3Gq
b4WwJe3VjsSORa0uUEc87zcPOyfU0p24rowdt8OJQtIoXVehSWOwaqaMtW7ONZpH
qnXor451pO+LiJ3N8MrUykSIBCZsBve/Nmr1jVX6mZ++YdtFqgFVuUGGQE/7VbfD
KUJFdOmPRH0OKUD3bedlOcc4W/7A5yfP1TQV/9cWmQf6OTl97ZZ0j4dtd1h/LESA
xrgCIPq8r3f7snluxCDqRgDuQK2r7ajSKu4EChU7Oax6UugLp7shty9WnvQzQIkd
lzMlzFqr5+l4PMtZdy5LzJvCEhJGrH+m0ko0Vz9MN0LoYNXv+U7RqL+V8HYy7Iz0
6Z1S9e+fkNOLvASBUfVGQQ0wnqNBeh16nkZZTsxlLqFYM9uSXDNQ3T7ldQCOq21z
tDu3YfQyOHkhXVQaqkx1avlMLZdS6st2T/dhpQ5I5CtuupBKLCaPnxwjwtHW0nMl
oSz06mRGa3Y0Ypx2Fxm5XCKWLFgrPWmvunRP6H7k8TUHuvJpE7wZ58EJf+4Aa/sb
ReJMp4sKRqCZCL2rbZXxhq8VWNceEZMuYgdeR3jxh4FgB/P9GAKkkJfFR+g/aPCY
r1tsozUYfgnG1nFzP+bVrZBk6qpLCocs1XQh/1SakgO2wBiin+Yupd+wBPTILVU6
GTEYnwgxJeKTwYH+xpjkNopK5L2nVMBVJX0rBLMeyfQLUe4P2xqIEt5UpftE6/8x
xxCwoGnJk1SjhBGQ6n4j7BohYxTtFyKh+Yfr4tJfiTbNTYLqtpdp01MLen/TCMF6
ygaHLNhZLNWJNm99YgfGVpwccnVoddGB6ejRHk3Ix7sDBr5Mi9HCfsCnktyWWN1f
X7zSUjH7nBmSymwdZtmx+qHtPO1YgVeCFVrlEbnaS8HGMQjBv3lcAaVcWaxx2luh
8lQ57HdFLwe/OD7phNOXB+oXUjtgvAmtAHYF7q2i4yv3KYX5On7ihZWqQJ1IaDoP
+swRnxURhgn1bbZ78tTprGfLMYb/7Tv5sUy54ZvxQIajnlQLdq7iwYtMp44+Z0Rr
/CTkqvwbK5LQVs270WLMir6/d02mjP5/IBX594CReac/p9VEyzJIpDQebnJbPYfJ
QwwqqI9cPAAOa1UDBeGsQK68OI+H/vN1J/9jgxZSwYMDtfJwUBjoLGV5cRDj4x64
xKR/Up5hp1Ie8NFx1/qtg+3ksyEAGRe0S89eG1plN/lKH8ELFtc4Bor8GRnOo5kr
t8c9dVaBUAUMAiJxg+zsL88CIgMJFJ40kPCOeAErB+pgm1DzaBHRb/E8XoZz2i3I
yIpmvs04RmWleW94KISpL9GYNbVW5XceNxjdxi6iJebUMo1zTj6Sn1LLSvnbOLIC
aeia5C4krvrrVTXy+YZCYcomxEwWLz551ZjFRY0fn2lT6y0hRDvACc6TS0b7vsW3
OymJSNiUTqx41MOTpQ8v77q1r9BwYhyrUS2s4FiAJzaNHm4O2kaiHHHJus6cyXY3
Xl1MsSq/eG+Nq26f9xpPRcv2tKhYbCHGoNbIn6swiugKNuFSqXTNyDX56U+Mb0VR
5j3/2uA3uqINVP7Gu4J8AzAhgH6YDjUfLCwCoL990RGDPavOi6/B23KxvJHuU/X8
u4LRyOvZfR1w5ClcCfeIhrxORPnlZ6TzbWbyRfOv0aJDjyjX80w1f8clnEvO0F7M
ew5cfxMEnD2zGenZ2ZUcDUyqaubbpVonLkx68FGm/IYHHrV1s/l1ifCsO8qWvOY5
9lyEs/VgpcR/Hce0/5kXqtWPzRQwDfe8dwp5Nfv7ceQgsU20ncyLJGlt89kNSJcY
HWAW+APzRMgoZ1MkKKUwUljhuMEUtcRBgQqmr4RvkwT7oVdFf5MOY+OIVuawnlmP
KqOCXoVdIybNdtEijizFpOvrGt6TEoagpb4sJZvih8Al1Et9mEMqRA5nPBIROAG/
z0GLj4TJ7e6AaZHO7T2peykrDouPZ7ankKwlQhoIgBio9rt4lnXC6wcV+C/nTkVT
fX9gp8eL3TnfGHxteZVfdxyolBT62CRU0QZHOL9MOEUI+IsArhKtrJojICpeUhGI
pDyjB+OBkA1hiYvRTVRvBtxupr1/rW8GxgV5tclOn572z5P8szS7wYZe3mZTKtR9
UQRpm4S4ope09mBq3Gr0jYWmnig99EZBGthiyGl/8FgO8ZrppofUuvZulvMVG2Hj
S8NjR6tf/66ax3N8H4Px7gtHFfe/xDLtQCASpRvWKd9/Ixj/TjyrfboOqE30CZgF
8gqMFt+7hLn4UqWfJuCixCtOJ/umrxELoCMu605zrUD0IDKWKyN7h7FuRJWdciDP
nsPZxSDlQlVi503wj6wG+OMb5EdYa30WGyvxLKn0/iDXBbTZi7+J+T5jycHg/kKo
6jQaMKHlIjmD0EL7H3PothsaWGXk1sSB5e8JJSrd6hnHhbVxblqLZM0xznbmtEz8
kLpyp1Kz1+kvMStcixqhQPVy/8BiP2U28yOaxzhX6Vm9VcIwxzZODo9LHZrqm7Ps
4RE9wJ8jA0MzuQaIydeWqyekYbwOgQhJCg2nW4ijQ0RrYctI5KVgUS3kg8I0HHNl
Mi1CcSAPL8S9qNNtfH6oPgAx0dMdd6s7W+D3Q4CEpXmJgQsbFXf536F2wuoYXGo/
yCK6ZvKHP1o6jn3WquamvHwc+L0Q6aP7FGNXuC2zFt0hSYelHBABdQsfKX/CiP4g
hB9mxt8K0LUDQm3u5Sls81S93D1SsqEi5QGNhJr14cC1nGY4J3Jw61QLxHGsr++p
X06gWSdbQY4zYfTOE0xU1jfccCY3/Zn+3ttTENrQAjOg+gRXwZOQPOkHuIPCqsgL
FmV+RUkvgSSOQFnBkLlMg1QhXoTEQo97Io6WsimsII40aqtOGy8gGs2cn5/CQSa5
8/hwMyudOq80a62Cd4W+B38XcieLqffMKcfkk0jr6hF5xO3oooC5ULxTXRlFlP04
LuAq5EnqAkCbR26emP++r/0KF5IxLWiKqDj5gGoc25p4+VceP4ALUarSdDKKhzrB
MXAFFDERyZSPmxgIC5xMJiAQm0H9ljFCwILQ4gwTsVp7j3AVX72FP9JShZ8pC6sB
qr4/QMpmB99TKlakbvb7AdrufIDzy5TdedKo94BCLeaNjDuAor8qe/vmMJvJ0kvo
n5qJ3/KcM/xlLwuU0vW3HHDLsxwwB7wqoUz9TF07dThNEEaidnyYcIbBRKwIH7W4
6B1CYUYP8p3aa8xn/mUPyCN0Paa8XNVqFvOLkpmlwCOAdlJp/jINLJg9EloBSwFz
GFXhAY4Hql/3plWYNTpjOCXl4nJI9fnmwKNC4jFcBZhDU24EFP2YeLPSqaU6Q5Ki
siV31qyYss2HLCs18FXaLla1GjBbjtVzPNbMFooJCi0cv1IrErU9hFSR8e6YYuiV
VWrA9eSTNtAUZeR12vF3teIMGRi9ORJUr/lRDUmL/WqlddAU8RA4UjhuyIoib+Yc
2JzLxNNR12cdrL3rXjxjKeWT8opJzC4EH4mM6rBeJSKOZ416SXMC+VJnsYW7smtY
CZh7svnFDi2lKKdE1qNFxaNWEWudTkyhtHB0hzUb3Bgx+Wx13B/Bu40Hch1kf1at
d/Osi8valjI3X7GvnqT4bMMmmw6Rh7FkCwR4lC8ttAGwqljvPguC3HncTnePT3j1
xjb7bPEcEqz5W9FHBfkOVDAVBj2dGgk5Bsp+9llBJKXK76zxn81PWw41d/jtqvW7
4gjKAhx6cpXnUuFKkgAgT6KtSnHbqrPooi1H+0jlTkNFkCM40xvnZ+tWONKYpnmD
E2JuS2gX+56a+tGbozPAvW/uZPsnPfWdxCguJMi/VeqJJGbBdkECd8VM96XV6lCR
1/JdJWMd71zMBo4joax8+0B5BNb6UW9KaebnvZO5umSooly3x5DMpFqCi8zwN6jJ
QWMm5IYNEbMhd2aDHD8C7cHLY7hDkeOjOzu4OcAilaZxphtFpLNFsw9LFQqi1gnV
rXhIdNIIGk3j0sZUFOWMyMOdihXajVugNxGq5i6OhoRechX1PyiaqcPvS0xewoEo
WYT/XDM4qG+KRvEtXrRKfq0zt6bl3p4SsQeMszs+txp5StRk2+xDvA9sY65WWjGy
ec7Ougw87JNfV6Az9juyoTstjTzdL1MB0Na+vaPA7E1cnR5UW95Jf0Fe1uLu69fL
342NZnIV+JAUw68sUx0aYK57DJt2ZF6+376GbhVCOhrtPfhuHzbrl+rnTC7q/lgn
KaJ7MO6oo+Ux6EhjfRPByqLgm6m190nKI6NwvL1P5WYXk5U4ZA/20YlneqqbeDAa
ZisoCnyGka2579qR/DJ/OfP7qBsErFQtkugCYGer5lHhgkjU5ZkesKdiTZjtyC6y
LmqfZOvxLm4j3JYF5sspwKGIqmAycsBp5A0d3agkkvSicNM/5OxpXybwhterm/kE
9t2HYCEKRTHgGXJj9TIRPT4ZTb4xeimRA7xsXDlhp0/qIvkBSHKcm81Ftez5cXPH
6K7Cn2c+bJg9Ye/+Tfp+Sodhydlak3XPeKQezG77Kh4USJYJxPTBqetciBNSmFPi
PaXtlDshBPxa3lZ+P1joMStrYAhuOlIKE0792VH/IhL7e68Chn84Ez+nUWCcMM+z
CcgGBq3WmGFu6rhS8+fSj7swCO+oeu9A2Qgtpp4aq4uJNOH06EX0nLt+Z1DyZQ7r
R42nU7wpHIs/DwNyczvNhjoiOQYGbRtQz+wXRI0TW8imXm44ZkHgPsu/VidwvDKe
BS5bNSaiQGdg36YyPhRGcbi+ECC5avX0/VliCWcAB+OPxyK3z8X2fcj5nxbXfq29
k//ulL/PxfXc5a0xqbukF759fMD6b4NJHmIPBM7ItTfct6QzHrVI4KPYvcqKAV1l
CiCp8TjjWyDd4XHXIX8S6LPy5B102cdKK3kFZo/MIwuLa1Nv4MlCHCa0PQTgghei
GY6jv8GR+zJBCe+KV4YOOOvj4Ag2z8QPEsXoN+82wsGALfoDPlqRAtfuliyE/BVX
NdlmL9tEkU6tMNnvAfrCcozuL4rrUf8zI+BJ0DamGkCR9tslE3Q+y/RGdfghSmdF
kg88Y5TduwIPCFWN8AYG8TqWuo0VFUljEbJofkiU7gc6f4yh1k8TRUVwnciFMprU
1dXebEYVMxGhuhI242VOid1wpXhlBv8nuEhJZCmswjUxLscr4k6j72JPkTS2Bp9v
AVmHjkIrQVuj78X1o8IB116B4cTdZQFmcMzDjl4UNuRm4s/YZiW4oTTqtP6vTV4U
rN96uxfeIogUbxxCsqCe5YGKsSp/lKQWP9ZerTFgAcRNJLfB+vEh26xDSU37iEpl
T4Zq+twdDWyfNcPs3dJqm8Sy3S0ffcEGXy6eGzHitqyNqFiXU8NR2h6HZDcRc3mq
EWL7kPQarqqpMltajjEzbE0xnEjP1OxJt1OJLSsTz5lxK7znzvprXBOrE/e7MJYh
uZ2xicJYgmw4RQE1qZCmHu8jM254wfDGh60kIWWZ9mjT7+DSB0XtFZJobPdmv4S5
SNnh50VkuLRESvoqlZDSulaOjaL630UzILoODvz4lMA9qXurrGoBqsul1HBk7kKx
4LFKlwoT4ceg7EpMznbYsQTxZk5Kadzp8ADpJltu0waXIgbFi1SrslrsoDuEzbVa
iqoR5FAle5aHDDSiJuJH50mLIQ7W0Gun12EFTR2/4BYE7kNsE8kl37qFhP64e362
LPaDC4tM6wsBrDAaO7pkV5NWXSzBIHaGHoSu8yqun6LwonXG6Ub2W487THK+U17c
lHeszyG2mDPA5SEkMzvbAtfohUZwDY7idmpROFPEHDYz+1D8ClDvUpXo3wLhQ2lW
iNJ5ktl7w1nzGZHCwEC/4/QV6C4CYauuFXG2i1xm4maU2CqY7PFsglRJaZWSqRVY
EN+/CkK8sQ4y6W2ToLAC1X9TkI1niZ0Mz3o36cLJI4syAcRPZQFJANJMezLT3yE/
L6GBYA+oVPSjGV6tnxzDOF8qszoldJJVTKxXU8NTTnkVJ2fsvGw3andt6lWKHxi/
JmCkzEyWkoT+ihc2vbnBAwyM5zNPoMml0xD84XXEdJ2grpliqV0wxaz5otTLT1El
Gv88ifKvTnigRamdVV0d7FI1VSj7ObtvnbuGT471NjsYtflteamW4U8Y3GcYbeuP
jRBMq1mqPA/pys0Ht3mMib30dxZfiphiVPkAB6cu7KKTOi2vRYx7UpBElqAoff+S
8U/53cJ1bqu1urXpVeU+leIsW7y9sAnVlMomD6uU2RKiRdmFQk7yeMcrvVX6GbQt
gJUycDX/3ChKmAftY+Z/ADo7SwkNTS5RL1EQnMY41FmguQ4pAWshaxXxwTwCj4k1
o4YVA6rvslCyaxKxi52Oy4SvGAsXpiH0lM37LCTkXY0Zt6yG5tpP5U4z8NwgAVnG
wUKB5rx67yJluAQR9Bd7MzmwZPfsqbVrBmfwUldd4GA8gp6WJy5267dQdkqMd+a6
8/cFc1ItHtjZS1zrI74mYIy2/LyVrgTQMi1qdEO2ly1JahHwYvxcjyBa6yR5OZTI
wOm5qlG1yOtjPaD12PVz4yqDnBRk+p1SfxbydledWWw712K7ZhxLEfvdaLx9B4Id
WMoLJSWhhgXBi0ckwtId0XWS2TjuZSGk+EnaT6xccLVWXtNvsxiv7yhNyyp+MOsJ
fMujFUJkYmaZOlRG6hvxzoYRbzTQtPZ1pl1SH4laje5XFz0t5loUTH0yWdcuzY6z
pD0NRlvWqILRfET2J//kHalvmkErieP8oJ+tJLCMZvZWNufpwaejDqcbHLVeYXYb
zMGp7zHx9F0E4MZvJcOBZlHIMltjmat2ztslGHJiAOwcH4metFI4+s10pYCtYH5U
H6eutTdmbQ6kx9Kqdz9o7udHXBdpEXSB65CY3MV9oFvBERHVG+8Nst5/EtnWXOgI
cGtGOen0QkM74GJrFkxMSPUmdUL3wMadH2BHMnMGTdYTOHIpMxOTbTPyg1aX6DQG
QUvyCV84CLg9h99NiDH4VdIjcKX+Lp3zVTKguy/CeOMbdelcsf3SMRkdzoGk377w
`pragma protect end_protected
