// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:01 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cP1Tm88ivNh6zq+b0R9s2b99Hw8+NRiwA/ZnUAkaXXedrtezwa8sO8o2vXEgkUpv
8vz17iF6UsnD+JynZb3etYuzfDhIV6HO81sF00px788gMifmnub7pDp413wPvd5b
9iz3GcxOsnKeyCA3j/kwERHmP+j4aH2IxCrKkoHx5yM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28864)
sg/y9yrefKJzc2XZA+6XefvxHCWxZjOAe6rbDxJPWJ7v2j6BidBJg/zfiPHul9aZ
YpT3fxqIaAXJ3lw0J9Th4Mei1hwDqfzo46MMv+551L9jMhQm4qoT+Ng42iBp4BIx
P7Xaz8RMRZ73Lo6wsLz0WG5iELEtHuk+A/tBJJj1mVTVQ0ePOnyfU3i75j+q555f
3pBwKfsjUeMmEi3Yf0m04Yiq0ucrudSBs1dwoyq4FnC+i4imNiClzQqtEJjVypHY
yiR57KWJJ+lNdfZYBWs2nRG9TXxkbT0a3OFmPEquGAI3PIw3i6UFFj5i0hfkQ/eF
JH4Qhm63NVMkMnliFFf1xagrF79OlOnWUgeYBfAzeyG3R3UKddjJpSV4JddvaqA6
ftMFgL6uo6CkiuN08RPPyuwNquCC8wLWXTvK6yqaMa5rPl1KVneCsj3yF+Gc53Hf
IUy/do5vaAyYReu5SKCk1U8e52wevnuiUUeL3aR6rdoO7TFA789DYsmxo8wjSkkP
01KabNFOwBefREHV+82zN75i9t3/ypWoKWU3Q7+LPtBblPlOGYmVzwqqMoLYkYr3
ub7W9jtFlD04uGyY4fDGMzXmKy0avu113OHk0hvalsVUvBgNyoOFTJNc5YDQIRKw
G1cgv9VjYQhcc1l3PupSfUo3wxsOXGGwKkCBgxMO4cUdrEUQDUmCBqMyhewWVQPU
ss3yNcO0A9BpI7noNG+gQFzFx3IXyreRdBJZ7GDXeBzGmC9bgK/5zVBQLdre6pNL
+H/sfoeRXZ0XlWKy92HPxpbBEK3QFD0lRtauQQJ1zsEgo2Y58uNaJfT7L6G+lwTs
pxn96cKgROx+yabuAgVH3eGTMkPXiTk59ItVAC2L8Xm5ISyCjDKyjAVDqq0LoGuO
XVK7PwSebH+ZerwQADz8DcVCmUFQ1ek8ICz3nUuT1WWt56BGrDFVOlxpFLUFVY9P
dqQRcSSVAnJtZUP9/p7FAW8g+re4l5tmAbzK0TzEYsiZeFcgdTXdXfwhlN0ShHHp
7KySeIt0xvcclsaavazu6dEJCwvBbYdsLS3l5IyzGk76zacf+H3njvJ+i4lUBuFU
+86wvGYLfEvnVpNgMjBtSs9smAnXMlTb+sQpwqv4k3nfcR0bMYYygt6xNjr4llYo
1vH/ZsRVqbfZvQSgWIZIhBZ81LdPnKEaRtt7UbzHT9cC/a3lqBf7Uv93BfYSc75a
uHD8jVqLc0AGm8Of5EW86u6cSbRYu9LugcHJ3Z5b2923og5WVu7ysnGssYLTbr9e
W47YLbWzTdWyZnLGgd489Z0D3KOe3AOj0danXu16F10P7f6cKzNnv4x4mRROvaOM
Zr0moIjAKqQ8WJnzEUrnAC0Vzc99yZyIoP9VuTwWaax8tPmn1Ko1ZcuV2zgITB/v
hemIhwm2Cpzi5RjQ2NMPt4m51Z49t1rPbWruOtsZ9iTFwf7VGCYKS+7OYbNdN+Eu
Lo5xrE3/akQ+yC4qy/Ufk3+EdQlbwMayCgvE39xKXiJJlofJncCu36PdHycIc3Xt
9as0qdViPeSGrpbVTR61Y9hT4V/pBZkHxXOGbDoFBScPKuDXhSQfkvJWIfCgNmkV
er9TjgvdjyriYyKNdiK1LxujQwnQWpiCIdVxV9vgB1bpqohkWQ3CyAvFaHji+UqY
BlH5UayJuU5EguYYi4lx9MbmVreRaDC/Cv138wZFkYpLEo0+ryh2bSA6hv5ciAJs
NP1Jn8UwKr5FxY1cm6xx92Y3WJ38avvfxTFB4S9axR6ob2hNmk81t2WGmrRPcPOX
qNupyvwlNJ6pnJ6ZYgBIn4UjyVqcNGwWoCIuwNWHTzUmIS2Kk3po1Tb2Owz/Bhih
U8KDSbaxh1bMcFS3PPd3c14nMvTvSkr0EqIZY8b9aNfbrndXgkg1ojYtT1dke0mb
HzhXv9fgsBub8qdf4a1mr+zVKIeurlCo8OEPWGFgDk8oiLNiN0v1aZZe6dnS9ftz
5gT9mBJ2P4t1GdA3gQ6RP0R3fPpenIioCrmPMHdl3li/KDgcmTtAyrn9S2MxEnxz
Y6EQi4yEi4Zsa2n5pMnBGjB37t40wtQfb2F4tyjJIVGPS2tqDtK5bwz5VUomQRHI
8Gw6wfpI4vtsHCqz0OLXRp20UMWNOAu6QSFWqUN1v8MaPg1Okqc/hav2n6ccdrvh
b/jV+BlsRMJleFbl4vN5FFcvHSBv6eYd4xvYxHAadmhb2pnS/YIPmIMLM4ePEtwS
QVZJrDeYKeBVTltR2gw2YtqBSrQzExZtiRzyRWckDM+bUYc4KYLuiJ2jLGFNGSxx
B8T+CryQLahDA+XCjrssmBPgtBPRSk5ozZI3NTiDI1KMXV12zsPS+QgIqtdHDhow
dQoK/oTHg51khamoYAjlFhlWRT9PdV2zpTFD83wtKYnIlG+mY96IvDOpenXXLUoC
XBUjxuyFtdFhHHhcFTXZheKaiJB8ymhHGeSBVkdA19BOz6v0dKxesut/iqzH9RjP
T5aGwlskcMIVHIyOFDsLU6UPgdAJAioEARdA947IsarnJlNuCFErm6gXQnVMYJFa
WVU+e6L/hmwTMwsEZ3GVgX1pT7ajPubdW0mqTJ9bABgJ1ywhkmOMKuTwXpllS7nV
+kpDJnpYITQHfxnynuseg/8ho0uiUVh+TKfU7m/ea/KjtXmLDTxtyf6Z61SZ8EMy
4uBW4jiOtC6r9CrsB0JQBooaVpHBOyfssm3j4BYpaStUhm1vamhVvKtaaSY5wkaC
+m2wC35dBrjo/1flHK/pbF5v/+tcgy8Pmn7+zf4kwpMeUlVtuD96Qe7q07RnHWTq
TdaZwuWPVqziG9VbRroxACQfDBDY75ArZwClDiSADv/DPZBQ8Zqwc0kp7YIZGQvw
vjdEjaB8Y2f5O/UIeHC7Uu34158xyS1FjHTwmS2eNZPfG/+3equsdcemBZEjuf0X
nrsyu7zd/BPe9LawEuHXLPSb1cEuslNTw7tER2H54gedNCWqm3NP+OKWS1TORCCH
WB+2AubMRi3MTH/NH/uysNwZigDVBg6LHTXPrmQ6Th8Rbzli07vIbxQX/iL6OocW
lwYnkND1AM5MN9+l+K67YP64blxhiQ3WAUGgHFSd04MjRCIK4TDJ4oQyym8vJnjg
pNsxo8oPW2s+Ud4cfBQ+T9qFLtAikj4WpNPSpv3S3P5+pcT7w+1iJLJhUVMHYsgA
kZsOetQTuGXymyWEb5QBZzWXSrse8zixLw5hC6gjAeF4FGcy9rTRTrYbWAq4nxDh
QUe2q8UzTkZCUX02MHG/QYg6ngtPg0Vte58lQh8NDnV/XU1pSPEmJzpu9fqmmJPp
FuD4xAS0boH/S33AUam1FT8sch7RJO4qHNujeWQynoQEbiOCy5UEy6DFlHcwLEsY
GEp9OmDOLMKI30yK66ksuoAghC0bJ0m26mMB+nA0KmtFVK9NBw8qtSOg4gWhov4M
sYNldVFBWTiWSJ10cKtS1gkQXXhMOBEhVFvXZRDZzFhL9+QKemNCheaqy7z9ozm8
RuzUMaWcjVOQYxUn+/NlhDAF2asKc6E901KvK2JH7E9U2vOBEfrhIPFv9y/0Gpxc
RXx29jYNBEtvHE19lleGJgVS+cvIsyIvF7/3nkX9HoZQe0wEyDabG+1bGbQTA4/o
e2oDnVu6+q365rWGJe+06jvM6BqOXo7SSsEDtKYiqGDGMvNNV0v3RiLK4bvuZnJJ
5PbKaoZobDgUzmZhaA9MQHpgFKx4JcfYUeWqfqbx62HPtre9RHYWUqK9UvscQ0eZ
HU97s7dTBHxQjhEx92PXsbPAJbXgzuxlej72xXCzpIYSbuAt+b9MpW417Mbj3GMR
HY4luEigTaYZG85wd2Cumh0nSXyVgA+NSk5ST+Q8VLsIWAKliSjMuY01iH/iYbrV
JBoauS6mRLnpWLpqfXttSGOeUc+HtG08tzaXzWSoZtyyWNwmxrZ2bSm+RmRKuZnD
Qmj7DeANT/WvfpswAOkFl/12V2uEmvKlFu6rvmGR1oD9f13z6Sfgo3O+XSy/XEae
7rl3GnXIv8ScUneNYTcdNCCa5XOlOjCKulQnZML4sQz0Az1cgGiR/qb6Yd8TIFqK
yLrt/7StjzPTRis9WeG4kzRNiU6tpXE4NZNyWWGY2DPH/UlVEPrxvxURtf+6uo64
hNpwNDehFOcf49DQ1xNk43Wy0kE48vFOFVnSzOkCy1bavb9+Ht2tsxZX8uWp6fv5
dhEDUPQ11SM8hOd6SP/Z+ao+Q2RdqKb5iX9Ks+HW+cPzUW7/IEkL9p5QpWILlwdJ
UV4LBjLitM7axUW2XXmFX6ca3FI40W/zmKzrG9jtecIMB7kPKLYSWcw39Hmfthbk
l4Wn1NFDafbySGEoet7c/3DGoFkRW/IHeWhaRktbqgAl5tol5ocYReIth3X+LU4k
LoC3BVnVdoHeW8uW3pyVmgZhxLrlZZoInG02Xk5nrAG5MHPL79bnaWo8M6hgXfRo
GauLHQUTdhddw41AaAnQsbcYyD92yJrbMZC6M2IIhGwv1ELnHDdsm8PoIw1q2T+P
mB3PPCwu4xGxyc8IHo+HEAuiBdTop15YrPWv24e/F4/N2UBqTQnBh9v17q8s1ZC8
HNEeatomzKL1I5x3YYS/Lri2DbN7fwShFPPA37MKNsGI1SjpS/WKf+JoPk6Tr+D4
fK9DE/8AeT5IiuNP6kykfba/x1HeAi1/rHNoD/t4+luS5NUnFZ3iCsi5gw5YmpbZ
9Z94Lr7yELR5rtglixPmgYBmsBbhkKiusWJbXbe+H39Rty7Jyx5hXToOHfW/GERI
wMYhNMTjUcVTsdPdbkFG4DuL65DNC/KupR2nxYjExKfIiDQAQUyBL6SNQpz/6/+Z
d+ktNFmpTK7LkZ7dh0+oEbC8Af+AouKAb6LffwbAulkdgniK6ES8rhSqmTPbNo1X
by65+flTpOonFddNliftDDRRmCNy6XJTPvwvlX0J9h7nR5jmclqvhLeysJk9/NEb
2eXwLzUbvTnju9SJjvPP8JkGw26Wb4E7W7yXSj3zoYkKoyffaQykT/2RfQdJqNWK
hQfHXfDDVl6rNZAC2qSbz4TQtx2sAUsYO0rQtio9nxXylq0VQdgB3ZC9nQFJTBBq
W29d5N4ma7gxsBFEKHTsE5W8+zwh7gWOwR/+HKVMqNm1CnwhQeXUt3kDnGhvlPaK
0L4joLuCbehe8TVj7yeLFwb6vsqUch8qCfArGDdfYE+xQhQbQew2ectXzbza0b6u
A81/UskGRT3G71jp+2XJoF1d20pafmgHHa245iR78VS98XQp/3NPchFEu89E0Tim
B3JJFBtEW0cYPqE++99GvurUzVHGENNQMJOXc36iQDeUd0VIEsTIkv7eZwSDSYaZ
RfBmbkGLX6KQnA0/zy8Fxcu2mrpnGEcA5gdt/L2hV+V+XfIYz4YnBuvRfRmy6dBc
xo7xu59nfj9YuSHfUxInIvJg/1d8051ynrJ4mCzGIW9WresfNA/YNfVY2fXopuA9
gn766WqPUFjZxmykgJgcWZQl/Aogw9p5zBDOResSH7+fnCYsHZcw8um/ps8q2gDS
3skRf37Y9Oem/JWBXlcHrbSX68dIIM0d/6bwXvWxDhjP070aAIMRdORgrHGqN4MJ
F+xmx5pcuHDlqMAC83Dmrk3Ij91GWpQOl4Jy4aGC192vnqEcNoLXpVPQ10tZdzk1
Wl+eficw51PMw/2zdLc5F2IHeb9CevbUcrG0Eld5KTQQtp8iOao26KN7KXMzbIw1
gry5cNJNNijpv4ixbmek21nN75vPKNNKp3oVS+j6UyNuVttsG0TfxUda5glv7GhE
7r2SBTTm83DdWxTWlYkJdQo+zXRpfTNzpvEXbRrGLNMEYrVtyfuXdJPh9spYnDOP
MOvR6TWFTgg6HtmF4Rtz0s9N6oW9da6zakdtMuAuUgTyjf7Zb8v0YMeE+jRtVxVH
k1LreAxqIvwqRYHthGoSk8MHLIO+dYS+y604dHpKt1jectvt4myt4EXRhUboA8+T
9Nes1KpTox+gXvu7JMsmvioR6zQb+Y5+KJXD0H6CLM3Mue5w2HWxbzuWGuSJpxuL
0JrkvN/YETBqZCGHkDS9LAlYb6/YTyQtWQy+TqwSVfxtsaGXEGO6uiERSvYLqHt/
VLcG0JjNc5VlIkdzQi2zERVFzqaYMhZAzfeN4OL+dh8bv+WM4ve5Xlr1HbpjNDGL
Lz0mWe2NhCq120d7MFaNhU/gmtMGTT/C32KMDo3nkz6L4KckXFnriPEIlAhBYf/3
OMBZzXe3hRRriNWliUKkmHiLk/4wlQvj0BKdr0h2Qa5g2DoJyghgcO9+dn9nErFk
FxY2kOP7t7NW4owweLVASd+5JSKRxRDqy6YbolFCyUUpHgH3LhdJ7vn0ARNN0hOO
ct4V9y1WdJ8efgGTTT8xyns2eJ0ZaBBJeeXACRXyQKz8btH1EnhJ+CShgzPre4Vx
YQNjsh5llAhd2JZHX5pxXGer6Y5wdZlxx+z27geF4qh4A5tOx5+G+UszBPu5eCng
Ok6aFw+x/5r6EZVBhevFaGfwCWrUwndwEasJltjdQJhb5+72cw6D19qAisx1MBO8
VJXqaa2gIXqiFXNLQGSRQY+e4RiP1oqy7fgB/ZSc1Cpqfdh6ojnAczXIc1XPKymr
/xCJy8fXhXz01SOVc5G11ERSm6ipJhbji7sTsT/Bjp0ZWy0aJEBRsQBnSH1T3FWt
tGvS43Jydxhr/GnQV7c/ZBlG3Epsj3XKBD+g7K4H7TkcRhDacPfMaRinYONwHpro
A3aD0n7poecJr8VHGExmEpE/7EPm+oJsVu9hvaD9WW0XaU4pg7uFPr+2ZljFdcKV
dJZU90URdbtjJQgkc+W4KeyOD2hGxgmAozJ2NC2hNlQKFVYtkDTxBOV2kp7WaOz5
Z5U01fVmpHEXVnAx6s0q2hLGlvsYFn64l6FZAxvUJEGIpZ7ra/IfqtdvAJDvAViG
HZT+HZ2DR3kzhggYmQoAwAgvQmopydHB/+AM6O60FC2cpd8ubRGgCP0gfo1Vpw25
jY5EONZTCG49fK+Us3P297rpN14qRtiHkNoWliPgMkfYVj8QfXb96tyWGLTDI1cG
DcD7WfvCcN4kBzukvg6dUdrOdDAb6K4Ha/Pj1tRwm+Ht5puBQW1+BwppZP6fkBHp
F1pS2HPkgbFvJreh9EkF2Dn019hQ2v96cMgdZyAbLkYL35fHNgSxzUceG4CXXtRU
+Qb78VFcRTHVmBGKPe8PBzZmiQxyhe0aNk5OTxDVUbhxO98QMBImVdYxRLwDUEo1
jlcSsvuyPxjkEic5JKYXM7BjyKrvZHLMnxnI/byOoGU8eHwyyGYWAW3RWvUJtNWT
GaqEKZL5605RZTtkQbjzPxh0yKMuoPWtmXbpXSUVXSYUOZzkZAx0Yyno9XslIppH
kqnFFstlyXLzaViLdOavfXQsJidSk+bFUQatp6BU12tVbuAS6QSHkRk4qfN6ODJ1
RoWsLvE6q10w2XMbjpblbpdk7HwQWaFwcoVTxTZJSittIfjVgdeBW5BzK64q7DNR
Nj+zTXdPJXl0UiOO9+zhiyhOXxiXRrcrKKo+7HXq+mMB500CHOVFDBvGtN03Fw7K
G3KecVrM7PJtfXrWfG+0Q+aH4lrbqPSRsixgZh8p3uYOWngmWnS4VZLiHNsd3XtX
qjvtQX00JVgu72HgJhwgtcFkT9CxkLCBk+ZmIfQPw9ArMfp+UQHrbLctfc+GY3W1
YBOKkD/kNKTf7BnNU950PFy+AbHZV+5//A4OeMRMxW8zpbQDyDK3HPrDc8WauY29
El+M7pt/QYXDHBIo2/QFASNHWvh9Gq8mbXIBG/DetqkiwLeRLlNuiV49fJMeo6ql
WI/3DAH8wIP3OWR8SG6JJ9ngw4pQBPB/NzSQ2TccJsYIVfAvCkU1YOd7KGk2JRoQ
YptKW9yn/tmfNpU4vJCMIBIaJFJxeS1cQLs19O6vvITHwi0FU6urGJAAClPjBRx9
nX30XKGx51hqpFYbXoPXzRdfJcRz1U2FQbj3s1lugdtOevboNx/gLrPs9tLYHcaK
djTpJSkI5lpmOshALf8maNjvfGN2tyvhAXxXIjAjKKj/97lLkMT5omk5QVkIxzxl
oyPWkaIERgv1t746X/yQpEatCJaHaCa25qQ/sUTSbb92OwjQxgXzU5CKG9UZ9beq
ybGC7cuuobpQl3JzmaJEwkzwy9casDf3q7lXxmO1/kDGugW2+9j1JebjxTAojEfg
ocPIJqxIW48eyC2tBBz8wdk6gQZE8noNesboeNQXmvCo1Crg76v3uPFiMucmsGvr
+FhrhdzaZIF7sBpRphQCie+0SBXhHWPZ/nYV4yeruRPzvmiOX1wQAdH6EfhaY98O
KH6lxUa4BPMr7sybwR2yL54wAnjPZBR+wbr1VTJlUFgPzvA9b2qPn9ttwJlYc4uE
waptSST4bXv3LfJDEBJt35dMZ4FYq18JG7CHmLx58tUWHS0U8gouPkiYMPW0V9NP
ckAStrQC6dRq+CRneQYrOLsBdS4Xi7UnfsIW5SMNFyNRIfl7V1PJ/gZUT+og9eVy
ksuUdJThh/TOE1it0MNaLZBB8k2QGTJ/bn/3+ZC9jY74tFqvagTyfFcMvsjySm2L
Me245ixMlxfJlbnr/b/rLZKthgvj67s9qwcpKi+Rl4Zmlrj9kBHRWYNCchwyUYlP
2JEsE7VQuTuKhfY3qQDWyjc0YuPLBgTdXLpEmdFtauaQCHUXEX+wtzb72UUM67Ox
sbzI8Yq/H+A9gIFjJn0aEiR0JAFxu9NqzUNjIdPwtOjOcbZXMT23F7YHaMjt0RM2
7GXl62OohIm/ZOw6BJCFsftoicKyqjBD+Jt4/2/FBwODKcsPB9DZnjb1QIITSDN9
SLOnckB3J4mPSQSkKMws8WwI+CnSgKvJgeGlpWKVKFoR3ebgmgPF/DekGBpVMpWq
Hs2rhgl8WLfTQ0P7FJeSn+Sh6D76fD+V3xj6yja6+p5udd+rvN/DKeEY4ds4sRlr
fO9V4sLpUXVjepnoouXBpZVxrszTn7ASogG0W2jMd2ZP40cLVR/7DZTnj9dwgomg
VIMlrztG4/O8tfBSRk9QnBUKhw2ZjH43i5MmGCqH8X/eX7lVWHbp9zwuxUeUFtzq
Hgkgd1iiQ9v0Amyf+x8nvWIC9Qnsrha3ODKjbZCz/wyR1WQS3jsH+xqaTfCwPv3Q
OZMTtEJEs4o1GdfBTf5sxxS/OyKH7l7zylDUIr80gmprKdwBNeTkmS/dAmKKkOe0
OIgK81i9kgCIY8PzrBqblM21qAVr3OdsucVy3wWZkvHyo3hiCmOzBZ5OmL7TwRpr
+tKrK2gk0Yw4jhBx0+VPm7tSh7HaCiQSJp0xKjd586SCryrEs02kFu+ILCO20OcN
OA2/ptZQdXt+eHucog2OlS7EyO3o4aHsAHsECHQk7Bib+aUze2f2EsMNlfvXvaSd
llGqAmpvgwwRLZdEoGJ1H0BswhGAwN1NhtuA9WS58ewor2o08oeGlGWMf/SMkI9C
wfyXquPFQsDBkUTIRMxF9M002jZw8lohfDzAHorYipUEBs+DpYAUa4UYa7E+7STS
5FoCAJ2PuKVcVEKq1BjfArJOp6wClDPGsmt9xFT62JxpCR0dFJpv22R8tWM80wnQ
sPZNWD1XJPfyKlk8URAIfsiA2x/WjlELEU7Fj8rL+0PDjKhhBSSzF7+h2zPfx50z
cyBOTerFJhM/nTRm4Sixq3rqyly8EPzNIJwGdhnJU8sXjIWN9HBihrITnM33eSLo
4776sFnXNJ1K8GAr4nluMW/5uQVJ8siAj+WN/hmHS1k+5AoZ5JqKEjc+OMkdJMZx
3gunoX0tkR5yZDGB4IVGtLVFA1z2ghjsw2x07+ajlDcgtlU3/51bYS5O4Fw138x1
2m7UcmDKQH2qTY4BUDrdZhzbGCgDz8A3KpJQOCrXbcixdW5rKB1esziX8s/iNQOQ
9+jvWfEMalAjlJ8h9+4X/t/17H1sKJ7skAt6bF6zCf8rHccz33fmCqiwNtnJnkWn
XCb0aB8q0VKD7e335lvBkjx+NY+HcZJF0tdUtcV0G+/LY1Xtm67OsGfG1tXGZU/6
wtfiL6t/BI5ggJPr6PYZ9dXXIE0fGJEcq9B1l52q6tkz/GDdCcb3TP5l3x1KMeZL
TN1n7HkoI/V2J1Mc/A9HYfl49oGswc1BOT93LKDTNZA3nBucr4PPUTviO+Q7lm8C
/SWqZRpkQ+//ioKQqSvhT3TkWCzz8lYB/HtPHpeU1PPf5TWkICFvXlW3Oh8UGKJJ
Zrc5rxLYgRH4/2kLlTtyKDP0l5oaHT2wivHefWEwaHBWsBDQPVrzVfnYHcZiPztX
eogKzNGd+9On5odZ93UJ9T+OMkzPQv44bZosaLng+KoOmGY778bfLXwN6XMBt7wp
RZDCD5JFP0mVb9JEFyBAz158kBSD0g7jI+xKJaJJ3LTfO5g7XWDLqoqSvjBhgIL1
NsI8EPUOkIk1LuUQP59saeqt1iCrQ4ZhWqEcRNKp0K7b25XyAd76iKuzPsDavb+A
AGMIMDAYACDvOiKDbSaEzAhGaB7cBMY6ElzfqxT6w90m4MXWnl0Qd51xzVqe/idH
lgI+oEnfO47csIX7Gw1SYGeSEeSLgsVtkv5VNCts0sgHJNAfFHti/2O3A2k14DTv
i7rcmf57uqVbipBczlQOHGAfvaaGjLQ6GbEGTBw4KB5Q9c8xuHDuHoAepuhhiOec
KVTB3pFklDqJ6xYQ9OiHW8dNhY4xlEtEyp95GtllTDlevk8e+Cg9py1jUZOBGFit
bvjK+91MpcMcKHxYS9IJ+902vI4s6w86TWF5RSUOARsMstSU/bI4cOgqJcVSXfw5
c4zGXBTNezOWcY+uC1W/cSrHBtVBTjm24XXWXvIjvg+dJnXWlcsVxmBuTniZ14HB
m7zXQp+sBcJMYMyCq/zdvzuh7TIPjGpYZ8H/0rZh60sa6xyFtV6COKrSeevkKWa3
5DredzJ7ixvuq6iqnaUUy9QmJeOTkJBwB83Cn0/Ulq8YhZbbnwrjddppFhvr74R1
a/l2l+9IDRS/7dGxEETcJ0Q+ZPtV0zRe0CkDcxn/nWSovREsUoyfU5hLZyvFMN4r
Tee5skSaZ8qWHE2vybXpmQYGOpdO9gDwtlD1q7IrmmmGlxmfNbFTVsx15tulDzHH
e0dKRI0U8nRrzpa0OVRYpfb+9/QUfRR3I4A331hO8P4MzmWJn0/qoK4onS0R8K7L
lxQs3ZFcVDSsPtyN09w9rnrFjUdm4tHihJ9+hfECXLyZmXOxBDoln2PXJxMvV25V
D9lvqteojNFBFPkD1/IgapyBxmH8yAOgkbM2aK+0zbf4n/kH7CCuX9SftauQjY6I
cby40BPngPPU9un8xu79GdGCi9i0s4vmcg+tNxA/r1Ysebf85tR9AYnQ3bwyejJ4
/1B43I1VhzNxgQkV8xK9SflCkdtVKN7g4HKjCLGGWjoXvXMEr//fhjCZtXdg2KZg
r7Ua/eASkTFVjdMvrRZQze03Z3inA3P8sRIwIEGhF0BKSlZaD942f0VqReEqVlTw
yNBctOI/sOY2YCQKexy8qdTdik19Ur09iH3p2SG5iUkTc5f6WJ1/5+T5Ubfq6muV
s0Z4V7YBJRipZ7unDrmntb0XHoy/DLbTiwAhQZqf4DixZqGCJOsUmzcUyEaeiwRC
jfa4EaoapsGi5+2r7/wQXN8qWnT6m4oRdnj8Xdb8P52yYy2wL26bsIzNjPFB6tMG
hTX9zNUv9lSqe5vCtBb18fV83/MAnysA4+rBR0y6ShqiZEWRTaGqUSTFC2LW29Sa
v5RjgX6JAvNXLdFM+rTGFcpSKnJ+KBfGLLlz2gW9bnfRKHVXrJEh9cvvJZYCLSs+
x/+2cEVXa48VkDHJ38UGaSSkdoelBOFOtO+RS0pLAQBJN95T0H7mCu0Zu+E69w1o
QFKevS1XZrtYWCCJtPKIGODIgj9/jz0K8Kuy9zlKLaVAH4AwPaBNwGyLof2jNN1N
jITRzXaj5+hp2kh+KAw6qnBlmuo9n/TsmaeVwB2W1YAvgjlrcTA39sZ/PBEpNRW3
jIeIOIDDNQGTF0WOxUNF4xUvBv/FVOL1Tpdpj7c5u+5jwk4qzdZXfUWSU5IEZeU5
fdE6uQthLmEhfnIKYfbgh7goPZpZWi4N6JaJ3Mlc7gCi6OfQKc6OoNpXUK9Geiyi
ML1H+kJSZ3FQnvcnmHnRfFUzMhc2AFZuX4wpHi8tgyqrmOKCaW7ztmGhDYfrmqlV
kYE5HBqDZzNsyK5puKlVELaj/4yG+jIVoOs6jHHcMPPR3dKo1i9mNVr9lnAWofHm
TintrV0SrRLEAlyZI5HQ13OTKiFk8L0Vg7FkI9noBAmFwfY9NFFjZIvZ8SB7ci11
Gw9e/TN7R3AKiNJpx+nyPCCDeIFs+WU4rSIVCOJppqDWfOEYCsEsh3mJ3LKxAOq4
TYC2ebAk4jEq9P0eXjs8gxc+DAsuqPwAYe08ydN7ZNv/9mcRFt4/XgNSS2b3fleP
Q+EDYX5fugN7HRn/Npy+MZ4GwLZEVbOi4EeF+wxrsS3RIsEfYG+biDunQuFWdSGc
1baecdZH4s4TaH/PeT6iVvYMYnd3dJdhgHBT+hlGO12DDAeMptkD2cHnvJsNIStB
kxdAnH7J5K0CqlGLhX6KNIudx+8tKPmxQyrhz9h/qBLnsFrAs9r6TAdx8GsSvTH8
rvd1SSCMWr9aebrklcJYwyTq0nEqNQDPI4SUNuchpfT3fwWoyMPJ0SIZ7OogHwPA
yhbVj7e+IZwQIK4/0ejepxeuBynYWPL7ccZ3fNWA0mLdbUZUqJ3pHEoTFtc7TfEb
/55kCISzZ6sxcRdTVR4Xf31WhU0G5oDAB+uMAp3Lr9T/RNxQb4MWb6tGxeA04Di8
rSHi8FB/f8BVQT68e21rQqGul9gd3DccMiwkc20W4dFmtsSi62BRGlLeXPXDgM8a
8R+Dkv/CWHWMk8xr869/cUpfw/ddOAo7SuTTD3yB09BklOPFUw/sCAa8oS5cVU8Z
KnhR9jKhls/aLfEO9Kod/UWHGiKhn65sQ6ICaoh/WFvk4eHlsk5VfUTiBMIxDZox
KBm+CVxJiVl2aQLqVny4LPTF+5RPZorYUufvBrd9tNqUdYPrDRUiTG+/n4cdjp1f
D1DhyULnhMg9tQDU4BpedB8L9IbCFaO3ZN7Ym+94T31IThe2d2YgEw55Tx7GC7F4
eM0jPvcgjC2vGFKOv1brnHPh4Mt9Q+C3vcFwx1AbiIDIebDrgB3pur4rgYaLaCFr
XB3O+MSeDyOOlCDTreEihemTGWS8G/V2wBlAxODJbP+MHPN4+IRW4cyIUoFORvEx
hnd4JO0AeMe6LqPrk6Jvp9P9UYCNnxnP3Fui44xvFiVTagPABkjV5nUsn0/S2NtB
Fyt7Het+n44VZHUO3wLk/WZ0FRLDUXSts49dzbx0i17lVFm+PmqhdZiiUCQUCWMM
Xxws9h4G0MUV1+P41yqifiX5p2UMp61KrwtYzQWLEE52RyeGBiSAdSYZfO7FeIOq
pYxNu0LS0Lgvk5F93S/pk4ZChbonCmwbWnKNN7HhVhehppCPDvrvnBFZ/yNOSrfa
4u2mbDWRaIJ0oJ1hdz41l+BWeeV2iHwzWK7lfs4uDeaq19MyLY5HmQEuB2m5Us7K
a46aV5ITemJ/ah1JcD7y6CSaxd0EUua2RLi9jSum8ipcH1l4KV5sttriA/j0aOGF
zImrqiZBUPI7ijoHTH0a+flz/dHHe6e+iD6ZE8D+pSMhxS5PF/4HIBh0ANuQF2J9
/PbBVnDzk9/RN5OdfeUxoKynrlDXuaH9N1Km8apCAMWPRa3ihAre7PqYBiG+bo6H
JkUez09LaT0QvCrDcWyn+TB2or3gAJ14lZkDb3+Q/VPw49kpx+c0rlS5Rm6OpZzt
is1jetALmWR6pIvbo+ysOLPwzEts+bIL0x7lw7KaklUBt1a2zEOH8XbTW6blzALC
g9OsXb9/oWVfx9XxarqSxLBQSDjGPh3Rs49Xg3QmFxUJT/kKay24DCsIRKAQ4uZ4
SsfWhtmYxah3wFXz6zYDoyY8/qVlPLme3X6tsONU4BFUSMW0dvVQq2LmqdAA+57F
ukbJfvufyYexCyGzuJEdXurcUtqAYnUrrFzAjwuTpYuhDhM/7W//rj1gUklaBIqC
KZ/7ksauuLQFM1wpIMrtEuNt0fl1eY4elb1WsZSZkl9m9/ulbTsl+cSvthvR9Fhw
WBYRY9+xLxM+DffwxCjTVxltrugK8yH5AZ+NaOwbyMV3i/pa31OD88mU4bUgY4qD
CcH9GLqfwEJdEZ4/iXUJIWl1fwKQ5DmW+cYFtF+g/GvNWq9mUTq90oVszp9mirq6
t3fwio7s4NddNJew+se3hBhsjuNdi01BmN8dJqndLP/o1t7ycQDqYJ23EdfO22GV
bIqt57zE2dMN5ZDivf2JUIlDBdMFlM8eXHfsLEBh+WM05Kz1zYaqGlCP4rZ3+Ot8
iQEsKzhy9dcvsDskVpcjigJYZ+4auzmVG9v13TSSak2762IWlUlT2GKtsshkYMiD
wwbl66i4pYdUwA2FiT5C1dBsELHAWuvxUg8PuUO2YrwOG+g2L89RJb3Sz3Dyk2K9
JeMnuk4W9ISJyyJY46XTZtLDNpI2iXkrDn2n75/kWUcWyMFhkFVbvh3Mo6qxL26D
tD1HGr3XiSIsNgbS+zpY6e2d2UNoiN0eMHOs5lWH/hCKYZE/iG0c0cs/OOopPpMY
7QMkcaU6vHJMvB9OOwdM5OJApSwKk1ckynQ3xo9QXLNwy2+pLki+ZTn9yTrIBVPT
JHGQKyrOiRsx0SIA5zVF/7GyiO156PCsXMCJ9W0bN/ztsOl64DoTK+xeVsxkNm6U
7REge6DZnYs/HYxmoFrGGW3A/nyCr2FyJyI8X8F0gS8N4OC5pzvKwcQ4RHl+ccWt
DVuINdlrVlPBylHqxKiGqc9EruhMvjKH5w77S0mXxeAisw4P6a7ioOzlc53K52Jw
P/tR13HaJwLDrPn34kc7qzEooTLIE/UpHs8/VllZSjFUh+v7TR+wd/oOANK245yK
AEKwZUsqVeIXYO8sU6siT4FED6Q78wqtVh9JZVkjCNs/Mk3bjWgOWfbBe0AUecDn
WXVDYfGD+9sVmnYNTOrFO6GYalrYIquLzgb3iJ1i7r6VZYJH2ze4WMMJ2bXW3KKC
q4ZrRMqvmqG7YEwlWXRRbXBf/mXpKqCniwm0yaV4FI89oSYMBzYERFbim8y8gf4u
vaFlG28mue26o87e9vndvG0zflUNz+CNy1GMAIlgSx9cE6XOzvKCxjXownAVC2Om
D6uwFY76dxUE/yW6kp2pNp8qVHiA2wdULo0BuNxmHyi1XgWcRKeGlyMz1B/QyGGo
zg1176aOr8BcxIiCe7RI+qtZWAdRxhIN66PGfKl+5eyfv/6fTfGVne5xStTbJLTG
Yg7CXV4rR2bliTWEVKSAwPNBUnSHcT9qKEH/3RZsgq541+GAHks6sMsOTvt3k5hT
6WM0RE0r/p3ljYsxPX/QvCxwcpzPZKjapD5AYjuCCKDydDjpGWsUSkBURpmKLkOm
MGuzfwIb1m1YgsZSpr9d03aj5haFT2JClfxz9K4bVWJF3xxdtFqvibFU6bpUgSvz
35Fv3ZawFZ1Et99O/3tefWfpkaRmEkB8/JovMfBHFAg8pq7HHHWEbqfWOxtTWIvs
W+e1K5aJKFdP+EdZ7gKdKPF23R8o651dgm7PGsQgU9zEUB1VOQjfp4PBrikStOHY
+B7Pp/Kwzo1CJa45PJEKT2owCuij+YC0zwyc1SA6UdhYWApWlmbEh21f8QPZKHXi
MIzLjLqs6MzBCwA6BSc36XWHB3RB3/n/Ul6m6BUEsyifsFE+uhVysDjH1fEx6Mwr
BPcDH3hrrrkaUaAN58xUE4ruqx9NnXqNPdAA+oX+TcM8bK5849eL78dlGU6zOZPp
kOE44UjwOJVZiDa4anX6Y6NXmbwxMWY76iCpGtJl6KvROM8cu2dfTC0Ef1+5NNL6
+6dYHJOyj8yJFV+OvUxli0rcDkNnPE6XJCsypBEXNLony0NG/hkF3N5I9HQ/kp+c
5b2Q3J6LleJKoj0ccLbgTMx+Z53V/qnCaX+G9HAkRBZ2I58nluwvf9jMd/qlscsq
uQ7jkWi9WncDC4BvBaGUfdGMPchUQ2uA3OnP6Q/H1Gft45ol+lXrJQjnZtA/sEPj
+jabQgZ9v+WJvMgmDkAKos64r0Tdaf4AMNKkpdu4LO/DmRxOZPrfZqSAX+y0dOCm
tdeZawXf2mg5rTYFMA1Mt7GEwZXOW6UCc+VYso7Yan8C1BB0FxLt265ai3ayiNiW
Ec2GPM00khVbnmqf+EbzzBTq9YqGNr0qYQx2oECrRVVzZyD9j0Vd6uvoGqsjK43U
6RrBC9M2lQXsuDRjfT6hdr/qzoRrpWxTqMoZwU28oi0u1Q9rnFUG6zU+Oec6U1yM
tv0yAXjhFOKzWrI6SpGbF5SEi+rIl65pU3ppustsyitl/f0hFKEu9RYrE/PvV97C
u+NCoZ8d/edqdl8aJOmae07b89qPo9BD7juk//5sKtZUiyky0NwA5OS5byQkSToH
tNGSzTzYQ4p45AkPdMx900egCnFLSuRaKrEWB3vrf0Tr7KE1HTMxLKu6TZdFyR0U
w8xS5HJwcUqg/zLzxymsaIeh31b0u2/UC+KbRcBkDqDmvpHE7CXYAYtxB2NTn/8T
il1F42O9GV6H4FvwwyfvII08eE84vrYJQEsJPYYqZxUpM/aQkaeHKcXay4W06c+E
f1v2X5pIxIuavvBMCGCMtDLjwS7fUPEWzuAHwHeQx49NxxveF7KHoAJo8EOZ/Y1o
B3jGYIS8Ah7jpaIPT0BCrFU4m1j+zabagUQrHdJEzxSsHbirWTj9+xy3tLz+H3Np
uWe3X/XcCeM3j/iG2whRR5PpPtZ+7NIvBSBQYPsOdNyu9BSSTUxPbHHqnmxZ/69i
zislvo5wrSAd9EY8uaqki2GcWc6452rNInivqQ6ug72xhZ6M38cX0JI5l0Nb+yMM
fp9U+xP//zeVQ8z34WlqMSngMYKnBVzr7XDeYD+J9gIxZUbNVfJ39escBVO+vuu5
U1TgMIHPtKbNeReRFMiIh/gczZ6m/OgOvjiGkYBeMdTEHKAODinOUb3GTJeJcDGW
sJqz4eQ1b7BmC2b3ou6alxQAU+vS2SNct3UIb1xFWlM+lexbITlPyyV4X4ZY9B5K
vkP0lOE8P1E+cT14mNba3Ap+EybBuNKBr+ioJYtopsQgS53JGybEMhUuf31eGIIm
YeEA0zFkMvLwGsoiYC182y1QCxBFoBXiTHXFl0BJwgHvJU1g0tJp+M94bO6E261f
x/GckoPTtpoNrZx0q0DDFwDJBiJpGZ9qdz0y+Le27vGl68jiJsZbAqxpR5w/XDcs
V/wzGx+cqqeLUVcGAVDc50U246bFJN07ZxuHZFkxai/OahsBAXm85osGhe6MDz3r
luktPu1/peswwCO9dxOpv+cPtm/3DxunyZ1S1ivyIeqI0eOMJ55z/InwJ7JViW/J
u1fjdLj4wmOxIW2h2QmoYY3mTFNmYcVodEO8cJnaYTPcGfgMWoYb2F1VGkXQY2c4
9KzX4UsrX1MhtKXlO54G3Phk7KGVRhMdX/CH0xTk31wW7csWpDixR80h1LfiIHig
m5fY60bLhmHUXzSlXwO1eRNJLZIOYaxo2PA3jPqe4oTFJ5/o6Hc7C2nuuNI98zek
9JQT6nQzox5DGumSfAcN7ft9HoZqe0pb2ocABecVe3cuAyXp10HeRxVWdNQJC6Hs
LdbUuM4DpA5GEWBS66zGhSKM4AmBwBSbIa83BTNf+1EeYM99h0vDIWs9LEfe96ga
X3Si1qVsnGV6wIh1FjbW7ODmVtneV4jiIkYL6VZmY4aiUEdZHUYGGCAAz6Taul7T
e8zq9qKLDMy4klP8ylB03ZqbrwLOizJ2qDKNgCzUkz0I9Qop2QcSrU9WOolmZnSM
cRU9RPlM9S7pZ3uUIKKfcjiZmRn4iGhrHkaaHzhHUVOyGoInqTLEGdbC9QwDtrgx
nzAIHlpDtZoZ8sw5QHutTQXsn3YWTI2h6sg1V71uT9LpbZP088Ju2r4gZlgf02c6
1ATfmZP4pRJ+4bqY27V/ggAihlnRqB8BBXmFibF8V81Tg4fmEw2hqk+SEeVg+DYR
D7E9EccDzAkkSR6HiBsOHe+oAHFoC14l5/mDu0UhkID22s10ZUBhMbVq4Aov50Tw
+cXjHM/RDfVbAbHj0faOEVIzkRwYCZrskM9fj/OSRmvm0aJklOW/H3KgMpEaRv2u
FP3XB/KGO0xMnpqGRm9CAVDv9zXTdMc5cavfDlAh3CPIoJejDw5T6hYLcu9uP7kw
PdRTgcNTbIP+tx+U+6wL4OGOZOS/46MOlAhQyBx81kaS7bpHZ8YzCSRq8kH/QHJX
imKKiL5yeqXRTf1sayxSE8OhXL93nQDJgcAWU0TNqZoCaa/hn481BY6G2gQCWKmD
rkn6p4KlkO4fNbc9CwwKa+DLLJocJjs+Afikm0/chzbgWZbpNxjzNZv0KbIxz4sp
QRHZyESWkaino6dnDy+JH9DHXbKl7mQkOJ3J4Z5Ubs+9NcGXSqv7gOe3lj2ng0Ip
s6Rjbgrk9x3br2zVKiP7oN2Oz0jDT+PztbRcrL9iySWF5IM286u0Eob88mmqivyj
wqRjI+3NOnAKrB8UxeADP3FnoABM9mE1+jVIPFBRpU7SZmvtLJ5EAJLz96UctRiW
FF6+0r2cYyeU3OPJlMm377jNUhEN1h++hveYWd5JRl2S0s/z6TRPvg+UgaeVcyPz
UHvYjv42JuqJDZy7vU9Ji7B8imWMWUfowd3HlaAcQBozg2LhcjFTzhh+cHVLe72r
eryzaXO/QX8aJXSB4dyHx21unaCpdxKFkQuu4y601js9SKPOPTuwn80/VecJYOVA
jxe1tFbVjqzU4+8ttViKFXjG9zjA+WEz5W8aPi34tVPlyWrmw6gq8HHSEcDnyNH0
WGqw0tp4cvMhoKtb+9t/nUH4+qob7FISI//OptKIcDHhekwsTUFdT9RaBWHplh3Y
m9zIywGUnBuXggbROm+r1phn1NJ2FSRSz5nCvBuR4kkWZU7FG7Gvc7Ps82TZt3LI
sDaB/XCpptpAHJ89g5TlT3i9DgKJYLUS+yDjGieW0u6Ll0qni/AD8x5H9W6BPX+8
8B8yJmanI0XJxfizRt1yWxj9utakYUWd7GFxgxhNzm4ydpKNPn/nUut4xJn7F2OK
VDb1WrkeLfV2A9xbBR1V8W1SiwuKOu+eW8EpvB7bwAUrb5+Ns+IZeemc+GL9J6/5
ZUaqEQT1mk+eBhfzodTI/ZPYFyVlIruInnRthwKruI0OkV869mR1n1bGNObK72vt
CqfNF3Ga1EtK1tfGHShf8m99yaGGd4Ok801RdpQy+H9ZjIYltm9Zv8tYZlt2BpJW
04VujLcD5W4pLrwe6tGlgnOR47jnjkjKktEppceXfb1ky2Pm0OOdMXB8xCDOVuZR
iuD2vlsaMdIAMxl+KSxsNHLjmrxICatniWkbJPmuvMDXlL8aAIGmKSQD8rBzjkSP
o535v09OBA8zX3HyJx7OePL96TJFWMSeaQkwYHKDn24+hBEQIi1DpyCzLd/AY4At
1KZeuJMyDFkDlei7QFzEHwZa9lKIYl8Imt7ismBCq5pKxzRXRPipTKxBeXeDrvDQ
7TLio+XCNBpoOHK/qf6RWuBqVyqMvu51h02LHNyUIyw9Km2c7wFJevDfJ/Ygyv9d
0UZzSAc63ZrZM5kPJcy5i707bEFg9JohZIoEh5bpaxtZcGBO3ARtWXoHJ8/JeOvB
G2tYrA39KEpoyUSkZrMeSrB5wmomoxDAEWpplUjWgbPPCjIvwFUUw5jY/37e54gM
I6DwJyMOyiUi9711CY7eLfFPw2O+JInqVafbNY6gqcqhCOrj/7YbiOrM6QrodGhh
woSz2+D6Pb1GdhmU4kQmTwh+wUifmkqWyElnSBGrzC+swl1GpKi9B8+qAgw/6jkw
n7ccIvu/cVoXEv48EhhqRJ2iWwf+9kjTObRvSxpoysKJzZYerfyIZ24hfl7urORG
kXpSAIqeqenwjP13KTc37EHtk6iY0qkX15A8/efXDpg1TQEqBxPNdb1uEythU358
vHFby45hbfitZS8hjE/1R1wHE8Mi/USQUY3elnUx4+ZeBNaNhTtS6tvNAu7M2zCV
1DeLE+qCdd8k25DAk6H9b10GyVyu0fJxkmylHcA/MtrgTJdBbu95NAr9jYzjGLfI
fGK08i6Re7zSkA0IV89IXxKnBbayNdbfUskxa1GFBXGnZRttSwkz1J94A6npJ7Wj
iwOQdSbG/Ma+NIwhFlII0TsRTD1C9IrWhKt9iAVK7u8UJXo5vXqzQXPRlSkcvq9B
OnTOAbNIDi+mo7gbcOl9ikO/JmH171rGmoSvdzy60SJoCxGTzNDjhW1R9DmPEKZ7
vhuTG05jia02J9SMf14DhIQYOSq1jQSHFrLXXWOsN5rDNs2uulO41OmRw5B3NQ5E
By2WmCfe/RA98JDeqXJnqQz9+e5UMPqokjvaiWfSoaH2eBuJuXLkRtnRqKsn2Sqg
nkv9+/mXJ7y6OON4m0BJr5u+CpRS/dHhlvp9z+Kwpj0TUMKRKKhQZJ57ulwuzBLA
UtDvafbiXfE83HR4zrm3+PjkjVrRUyKW9Jp8EVFS68GhoQuR33FH2TnbNWmpB997
A5c9mSDHItaG6przTsvk9ikjIRl7oveveNKaHc2xVvaZRC2AX0RipXzQseK54WTf
ZI0VQGmlOgJZh7FAtNYhfBPVoBqHR4a2LmTHwK/AphQKjnd/t7OgcLQhC+aStuyu
tzFw9Aixav9AyeQpp8x0oUWCNMJtwujNMronpGEL85XuXSMYl4QgtKp6khmpEvn6
f8x9N1Q4fb7asmeMvf4u7eAMOdMSZkhK/M0hmwbxw2TU3UpA2uMjaLaBnvin78k7
OGF79rcpjlvTfvDDcdtwcaNx1T0Ub6qXTK6LQxHdvvGes95sM+S9Gn4dR4jR09MG
5lt9k+1XZJWEUaqHbmCWql3RvfJdhuIj8ffx7LEmvDHqr3kByv/78ExxakAjvHW8
UmsjC4ZRQ40aGDqv4kn9fseEYh2vkwvWLOH4HV1SpbYKEgwC+oAkTYExmccbCBLR
+MasLAVsOmk8u2Sul6gKBapoVoxtNRsdoFCGeru3/IKZA2tg3obn5YFxrHlg/ao4
HxrC/5uXspO1VgTpAb3HD/h43XG3YnIdP4nn7ABzMJkuOBzPDZxU7EjeRnoxFdzy
uFWR1yPj0vyIBA9avKWvJ+L7M9K777BbKGCGEX+nXnR6QHuykwsMHdZcKEcjMxXG
sg8lEtBAsVbXinflz8In24bwddRiiUgxDpZdnwoewTHytvvZYG8U8183uJgevMgL
yDErj11gM+cCT0Oe+HSwG4QVsvKOxar6/gPOtLoxXN2KvCsFtEmNed9fA5Wy78nl
kced/0J1GWFqS4jZNGGH64pPEMhlNK3SvrzOKOAz95XA999a3I2ImuBjfh3SfXif
5ZcRolcjWc5aPJgquM48HTKHJgJB1gHUnWCvEaLHY/ymYGOPgUO2CjkyoZWsQSWj
NHkmAv1vbmmHzN5FEqEwxbBwn2BXJqzPiCVy4vxD2kVl7EHjGEaF0SrxCHcJWjBp
ZSalgTBSHKw5RYydj4FegTi61j6mGXdSaETWPTSQSs3YJXGoHKl0Kc24zU4+R4MC
iZhNcmYmUQr+slRmJ+NGlJhVZc4CuKozlBS/0I7oj0PO/4bTms2qds6UbFJt5GCx
cKD3fBuJw6Ih4HepNgeNXO7zWX0Ijf5PQ4/V67p4hZesL5dGSgpVSYn3dcPjcv08
EDg407O2zBEhFNZq8ioPUQRJNrLU/Mfr8bXoVZ8cVpXrACCZ64ySJpovQxZ2psks
pc7DSOyTBSALQt4CZeUejTrJ7dGKwfPtEnjcN7IbiO/6ZhCTEHjM41F+PBrBZNra
pTJOVVejMpCHt7me0F+iVZDoTHe10vKKT8ry5uHT41tOM+LoHs12V23YvGzfMUyI
WU5hGqWTxJOf8ZJZT64I9wFktfnS0MrhBGLaNgqn6qdZUG1NbEX+9R3487zJWefg
N5oxQVwaL0XQlWzi+l9DayRgtl9+aZcvS2xzpg87JfR1OFL0hn326Pp+JDbM+2Fz
CgqWe8I3AmUhXCqt95x08jbb0BZhEogngvKA5edbUWa5VzTrS9CsEel4S2W0SDGf
xh8af+BeTql3WHwN/G8R7k0mSO63m8YPNyjtZto41Y3OWUI4N+3hChcP7s5ZvcFU
p48g3d+3wwTd+IMSRp0bPnpIcAsHXsujPRsc73TNhJbwGI5LxByVoXcuK+YtkBp1
1RniO3PQPeed0giCklFzenJju3VrMycwq50gMnMRULlcdIDtuAKxt6p/ZFSOWHJp
C/dvtxG5bCjYwOEczErY3QSFosnV4D55UirtKfaqv+o0Mf1F9kD2F2DNnf33USvu
/K/O3SlnaQIzdXk4CI5dpNPNbXFuhkfRwn9wLyCsSoa1b/YCqaieG7GKpzrNG1a6
WqA6pKEjgTPtHFXPniKi2dF+iWK7YeNCDPibcRlZTRQMtBApp0jv+2M+27z1PB0j
g4edS4H3ZRsycRHL+O9Zk50sKqBkopm70B2ebhH37hF4IqrAWROUHKQ6JScV//t7
Y97ZdVhUs29MiGEp9hqeyFM3qjVdYcvN6+CXq6A1AJj/yw4LsE7yZdby4uvShCwY
cQsWrnKz07jwGXq3UZFPL8GtEWQTJ0clyFFQtjnH3te0MiibToTSP5iwVSvebeMM
RPBQio56Av4AYmWqIM3/ns8o4mRZqDgFyUaqVuIWjbt/Q4V+0vLoTGvxuTWYQ7yy
PnDkBp1WPZ08v3gB35QQH0ecEsd4mv8Utpdn4deI2nudxxbhWogR/Y/GKwMhuubh
nwymnDmOzja/G04F2PHzL1rBguYMhj3bvDdM3bA3hMl4P9gsMv4Knj6Du6AGhBh8
ErcCNrL4LuphT9+7rEinKQvhQLDL/+ETx9nP3mKKt8ELo5QOGxfejwBhgG/2jEHo
zWWAP0qp0vYJF8lCjoK1HbHlsj5efhMSjlpEJoCB5fJdKPNLyZ1EBJZNt5TMjJK6
v/4IF7gpxjDMsSoBQsYu9cb+m5zMItfg3PxTx+EScP/DbIXfDtlN4LFHw9MtNh7L
pGranollVh1CVPp/SvoyC82PMms7vTM8u3z9eggAHwwQWFjbFmnuY1vYp9q1zuRs
5soKD2oSrjKVHw2V4wrW/X7R3/ILaA2w9a9n1ZA9Hf5mhckqAZw91Bm77Xv6Apm8
FDZ+sAOqTgyVKyxjgEEpFyECYjVeLHCNxuT+e6aHk7Z1Vf0VqJHjQr+P9nKg6RGQ
DKsEESqn1tt7HB1mbC69SoYDl0Ixk5OsxNnOQWQUOzhbHAW6Q+9jChqQtR5rXQ19
78p0Uc85Dyhg1iiw45M0OgHFn44B3G4myNfUqG0+0F0Ul7Vx1PLso4Rm6Bm4tW/p
FTvxAqbXyDO4yH6xqIF5FU7+Llzx5wsdYJif3i1OWCqoBzQVz1XMt7xsdVEjx5ln
Rgn99iuLGc9etvY/BQ2VdQHtGuRpQJwA2Avgb4QrgZkF3+on6ZvQCPwRM4P0fM+W
CzbMfOHaatbWx+BplO79P6tfAk4QUZ6aO6rn9sMW7EwM2a/iYapq/XPeJWe914bj
k5Rl9rE7KQW16/EahN3Y5AxK7v9rFvw51LmbrlpmDruYgCYTIGClJeZ6fqT97ss9
5Iy2urAYOPku5P2ZZZhmJJkQ7ym2armf2sBHjOQZZi1k+3DI4eG6zkv807lXaBZu
zNUcwn3WzGx7qzPEC2CZWxWiXXmd+DsdhFw9hR3qDw0KfsjFNrUkU2nb/Ba7MazT
aP4wet9yP4W4ssnEOt5/5HxFamIJnTR0sSLHP81+Ii6gXDyIWWWAl6rk/UDG7pQo
B7TngfEKE3IByHvDZNCktS1WU8ORE0gB+8aoJpPfPXg//KtKjdgXJVvgxDuxSh1T
8x+VEiRUjaqQJ96B/GxEJIRVrF1ESmQRjmZIa6XUi8NEgYuy6aJXkO2e/iUoPMI3
/YNXP0pLNWlEhHOcvZe2jZKVFHvki2La85NoQ8JyqzPUezz6Vvho9sRxKRTkOM24
nHLEZVC42s5YfY8z0nyhEn7nNe3DkSFeUSCGDEZeTBL8Z2zIDiRjhlSKmGDGuy6W
BMhzWD/bR/f+H+U+TgtDr+pDuDeUxnBnSYHQj8f0RN7MlTxHIDj9Sl45qi7ArOOh
23Ds0Arfc+83I15via0CWvSA7I0TCm09BLFTGuvDj7xUXVPhPD1OfNv3NyuxlUpe
Za/QbdacWn0JnMqAOoRBJUU6ustQ0ffpaQGuS7TudKZRvIvGmHrtZuO2r74NQ/qv
TI2M4oB79TIoW1uG8dNHy/ybSJPWKUs2nkMkeIpW3Ee1x8rEjiTvV+XchaWZtiNP
iJwFagHPBMWdWqP8C/mUucTpCRSCJpnEX7xVrBLSvcUMMqw8QJ0RUZFkkyOznNkh
g1Fvu00O0CN8/q5vd5MQUjnNJvEkzB3SDL+RbIYOreiEOZo+uFd8eKe6cqo6/ZNT
0Ft4xEKCAoiVaO5POlRbRUBnNdJzGWvTp5F8Y078ggmAZPvHbQ7z4k7548+ceppz
Tc6ME0RFa8nJBCoOMdU3qNVFcS6cXG2pgL4ifGhfWJjA0GjQOFgPmqOhe0euVxc8
lzlKzuQ17fXAolB/RKHgSYtrsSIc6AAfdgqFDA8gnbSD/qfB6ZhkR8heSiiVy1d8
QmjBRQZQKGmNyXapOEGKnwNhcJQ/I4SyYHHPrsv+VV//MUBaHxzFTwZJRxh2F5j9
zeSXrk/Bol5E+oLsxqiF/O52g9CM7Og4JlILxQdAy37sRMwJw8Fqp3BOZ8n6me+c
3ATUIZ0MzHEKIQY9IsXMkFKdrPRLlMOqg0koW9m3ATRByZLo4BopCcgmAF0c8/bM
bV2/dr+z90K0OAF838yoS4Chwq+p1duRqWfn5FwKndnXxMvWSgIeAJE6Q1QR00xW
edPf9Ftfv4bUwNR8knWU+TBcstKtMoW/3DUdNMAx5m5UHfVeNURVu9Io5BcXlsRw
ywxLs9/EnSVfubpap5RVWTPpAszaPCww2G3HyvScTwcvsQsU6KN7KVKADATk7RVG
iEzcuD/qskIM2J7xqBqmhf3RH6U5UGBO0w/3gBUkL49OZiKnNfZSdsLqs9Xsv+39
vogkkR3YJd8UbtRIRRSxHlIryCgOdv3LIPlEtkZkjyobRstwoUsHpBJAoFbZW4uc
Lz8KKbJgzblrkHHO0TyFuHTvpOWm4jpf8IW9l5D/owMryqlVolc2GfQgUvL2pD38
+S+7waMiBlGlSMn8maNSWq4E7UpoK+xS1MOrAtHK1sGEOIpF3hkAvpxOGRNjMVlM
5TAIOR6XHZCs5smiABxX90fM24Nolv62PQGsEuVKX0fGAkS3gxBLn6FoFcb5JMyH
7YdgJ5vhRZSYvnXjd5ljbB0DdXd0e8UCvLx8za7L/kD+8rRFnVpWM7MyCkdTeEeH
E4+t10MxNXPNciA6I8yGy/JBQDUm1Yr+P3kEdVQ7pps/8YtgnbxMJC/kYLAzmo4x
9omNYbb0xrMSIxUFHpN4lQDn0v54HwGEWrmJLDH33xqdYe4f/nEfaVndHsk8ZI1o
D27Hqzt3wu+4Lj7pksQEGrBwIO0jrCK3/fnbYTeuPO8Cn1T5/Rp5xPI5Ka25upF8
+cOkX09pjUrjDBswDZ4pZfO49ZmOxifAinIo59MfON4LMfJ+CXe40mXlyB0HEkgM
/vRVrpf14sycb6PDBSTo/lrDbjRORoCGvazxaaR9gBj1yQZhupl82urmjNF6S0dz
zM8GJNW2j5rYpGDpjKVWATKfAAIPlvJMw8dcL6rPTvYrKF6pa4ciAIgzXqBYJJIh
Zy+zEug7w+ZHXrEIUQ6Khx7NG/iwDhxV3vd8FuxoFgPlp6viFGVbT3t2mWKNZjBQ
J7iYr+JdprLQ54GPPrl39WPF9ULADl1EXFFwgzqH9FWO8sxOwzgMAIWrkKhsJfID
zloA/2Y0d0BGexXk8fXYq6sX12ceWXNkhxwmMMlDeCjDp4NnwPfJ6LfFkpNYRVF8
B2Iw5MS6Jjc/JD6FLJRgJVgwZTZvHg1Rl8pd0+aLaMNjn//7/VshAKMAw8nNGTcN
fBE3MXe9ZDsmt6nzEzzZNfDEBGqlZJSOI3zAzafRua54qIINsv1B9Kcaxjtag+ho
gmZADaE1EYoyOPOnrkw3So39zO/gM6VlkGE1c/DL2mdiZzynO5v/3AUqsQ3hX3zN
tlaxFtlgWJlanubK6mEfUMMidXiUdCH1p//9//bXWwel2rrDp36dhOEacVE8HBRO
epttZKba6QrJMzf5Bzkv8l/FrBrNmnOk+vxIr4QTLSLpJZDnR1urPR72fNdpDBa0
a9aW7oifugNzVmZs0Rb4/lE2E2UBiYgEa7X66gr7M961sOw7wiaC+X7vVjuuWerX
toij2QpwL8ttISL5mhQzRdCGHf1RJzaLK0RiyFGZiVa0QCC0gfUvFUauSBeXn8LH
ObNwugOOpD/yYGOZ6qd1HMnse809dJZfCITg171iJDtwwR8znEMrkmPCof3SNHka
RDnJ/CeejcAlGha0YHVxf3MAxBBSZDFNH90s7rvvEft141g4kQVDByPOU6ogBqKR
My1fsCM0IQ/WrdednLVa/J66G3jQAuB4SBJafSKtIO83zveKfkAagozQug/5rFmy
s/kRqTHvxH80lXbnAPV8swqn121KH+ksa5PzUwruVB+W4NrnAuZE/wnjatEAQ56P
KtVe4mRw7MkDnP0zcfw5x3UKhNsRUV69zQ50Ad0w+hhA/tP62YXexiP31MS+0njq
QSNlccW8SioZW6JxQOK0wKSOw7gbzket9485SLHIb+1MBiymhvOlhbDy6A4unxKP
/jJigIvNXyAOZQdFs7E48zSHYrIiluJju12RhCcdLjPlojmE83zGxId5TPuU9fCV
bIcX9L88u91329IImwTIYHNa6t/lPRsN9f6cR3F80B8LuVuJRoHjZzeuJmbgjYVa
1hWTQtYruK8FUH5zRXnRExseQzSYIiJkXLy45250IfgJ5X4ciZxsYEthtmz4WIzm
KZtHMRco71+cZHP2uORm2EbxyEU2ueaLw/GbBTH59k0tKuawzMC8G8OvhaeqxW47
MQBeCQ0JpztI6j75PHJXKJAOMyGCjjkvM1RqVJdyj+0wpkfExlhnxWt+Ned2+Q7t
p31wcKmejr7EuB39BdJ5zBrFb6E+LyexBnGVVBJTsGDTUoLGc4arBTv6NJ4pZsp1
g8eeMMW4Fo4Mvlxc/8ndNZ8DH8pbV9q/JLElWa6DEwbpYERkAF47YrdMSRx3JYaC
SRHiR/eDqwQFsJMzlOnKonaco8vPFgEy9id7uy7SUhWhv3Zin0QpKPtH3AVWqqFh
/3rLLtHLqZEHW9NNJ36YAr0c5buT5mkHUY9w/QZXnkvYxwV+49AbIwtZD79Qin5e
08Km9qWGrQunxQYbKVkpJH5JB9s6dvvVH1nVh13o1U8ks+QGlw1NJdIBNzsppnY7
xZ92EEvB1pS9oHxg4UDUvRw3vHaq6Xf0lLc8kEMfanJQoeQbVVu+W+MxvuUpQHLe
vRQi2RtWRX/lAF1dgBwPGV0816QiDJDxF1ajh3t2w/YCrsmX5d6yWhFP4W9vc0/X
yZfFqjQvH4hUxrQ5Gl1O7/ShwBbV864wJl30o1b5ifH4GFvaUmm8XfI3AMbWb4u2
tG7VvMeFilUbAEFZVX3xAKEd39tSVsJZvMwiC13fBKJlzasNrZ/CaEiAESXnw9/8
Vd75lSKBIxebqV6D5ZzKaxLhLP7qriBWxF34TVyT0MvXVizs6RNMdNeHBEUy7lfr
wUrfDmxSGV/4janlEkWGEfiVccV9pDOP9T5nVoPHUy2Me27Iln6Wb767i5aMPZUL
BTCrI2pK0Jmq8r8T7OGwDrltiin/2jhX2PDn5o6L2njYmaWydYy8pwmh95v8D/Nt
nsAUuV4k/1P8UfuZMg9l8hmpp+PIZbvyH2HX3vVWFroyM6QrbfU0BmY4b7EWBzfy
XgV9WaNANQVTdYmhTpX9vDT8HkcstBzFjVpg+qmFajei+U42MxuXxlrEfs/6lCoB
yF/T0AeQu0Zz2wibKQdCkppqWkmb/mJ1kPsEtnIh5eLFvA+SnTcEoS/mA1hRZE6d
uYW3KzFhrnMHh1uXlwNc2YZiIpZgsig+aNoZzpP7JPSlvXHzaNN4olB8wsi0qyLi
O6jK/gjDdCQ6MTg3q9ni1A5UD87j/8O4wstJxA6573se85c6Vdw6lH8AnULb0zEV
/VM10NPkRoa1gKuxJk2qnfAe4IIglUxZKJutOYoLpui0hNGhGpZsHs22OnXwor1S
pYOfCU3SItaNSdeYpEezNeE1yAyFnxNHObjipARzgcS2rojD02/EeI3KfMjGr1DG
vhaN31DXmOh5OHlGhlalOLDKQnW4tDzDH5UfPqUrshBRGtlihW0DDY4j7W+F3kvr
1VENw+NSkDIuTkVufW21ixi+iQrNRl+BkbHev5AgziHqkcgzcBN3hCAJb3tVPLmV
t9YdugSOjVk7b70gjlXaxv+tUY13EBZJDLVRxa8a/6fQbKlZ812ZXauUVgCijhzv
HoIef21b/O0SLTL5q1EbeLKv31MzK5FjovKz3iquvkcXpx3/7oDMzN7L/R9Y//4T
h3b1fN6thermlRcBYlnfK8+lVC78gi/GEJPPJevEmQifH/pTYMj4UxbNQeGaZKwc
IDlmF2+vq7yaObS80FUM5BmVcb05JebnGaLE7dDMswQiZuSw74x5mrYwT3JnjtOd
9G4bwvRhlRRgIn1Nqv7XtO1IekrwgrxF6bOZOenGUrHgM638xUL0/ZQDe946uo6z
76+pMyMuxiIKGRSVY9DF9YNN+X7GUQnm/WFcvEu5Wi1EphXFgMfv0a5Hr1OHq5JK
EhaLh2VB49Gti8Ou0to3wlnN4HEz6/CcAK2e8LV1JTN7Jws9ozu7sIqpvxGN1bMl
jWsrHpXRmshGfEMQ6v1BH4N9fiSgoijklcOyywiR8yMk8+hkVMNybLWZQ9vPMaD0
neEjdVZXD07rOQ2ewTnrPFQkJkjAkzKN4J0soIiG9e3HeK0bfrOao47lx5G6qZfI
+sa5AoaJRfMPQZ3iuo3cRSgmu59NBZj7pCCNZyocK90f/O9PrPiwHDBxAo9RDZuF
PI+QjWwSDIpqYbz8Hh8s1GBGdiVTnGC92C0XMIPgT5ov1bYKVMbNulTR4dnLm0J1
wd8rUtNUiu8Hh8PU1Zcr6Pne9kMajzi80LBKAxucGFOWm8zJ+fEa6rk3TBqeT4v3
OpxvhLnuH2jJK6tLW8jQaRmfKYh8QHcMG9j9KFvROTwgQ1kQ/bgJwyd+zpwgWeEI
+yHLkiwfIURHXx0jkLnU3bZqDmqS716IwQWRauFZsIqywkcDnNiaFzU3TBDzAmWK
FOI7r23y1PK+Qg5MrmJyIdXyu0ZJqDE/lTFitLIudhuEwwRuDrOaM5TQtWmpZPEj
jHrN6XeCd0L3qrUZIPYGQaEwv1X1cKepGjupN6Us1LLdBXEkJnxNsh1rzEB0trDg
j4/N77GJmMN/sAl4nTG/pUb1idD7g37T9YEEvOoD5onciqLu5VCuB+p9U/uf/eIw
I0PCHNRkxyGv79c50cir1DCWJ5FAXdvZabzA3btF7igzOYrEmb1VDPy6ULwuh2FQ
eMQLLeASSzAwnbxRGOIXmuIQ6NSnpH/4T26V0WbYn/1cC8hR191CmShFToFiALEO
dUZX14qRIgjateGx7EeW+x7UCN/jR00idRYXOIGNYqsflsD2xcai85L7qXldmbrK
NqUGvWmY1fsiM6vOWA+CBJbFz0jr/xUNK7EE1mbKi6+aA6S44I2l4zeIIrh8rVcF
yTRL2Kf4QfYdWjJ58gbVwPhLBx0WeBYc6IKadbPPGS+uJnQHMURGIIhcrjv/NnO1
nKbmMHOMS6p//HjIO+zd/Q9XDmipdraqJxLjED/nhub/e/WHfoE8AjhVA5DRAvhS
xbBohN+8unUaB162yk9gp5H4k9onuanXRm5H6e1YzgqP66a4NeuuAxS5obTwEpHQ
/iV3zOieg0YLRrx5qPCzNrb/2mfHtPpTYyb6vsPE/4fdC/dT/Y+dIQfQZqP9/EJu
6Dm8QFjEpsrT1VZdHi4fPzsubq5ocnMCSi+Rr94YUVDy68Iu2nM5suR3ZXZvoEHY
DaT24meLEiZONC3M8v4Udds89EjURpOe6eZJ+pFGjVmfBevB20sxuNNUlAGr0OgX
tUd+0pnlI2hSUs7JGz1pvkPIpxU8AFtH+UgGZJ3/Jg7ioa5NHOGgEh7QYV80uAR4
nCFJ3SExw9mdzoGuifm8tXZqx/Kya0/DpRs2ky//SMHcsPYSmEn+qrvJfKeamfPr
+Teb2WMwCmPxGfuUmeSkrpKAlRTwdjT0rsYttuvWMOGYUmaTRZ/rxB5+jo/vn93Z
kTX/pIaeEqu9bNqAESJRQ02oG+6H7gxYmtlMLLSTLp4PKSaO3khaA1wrJBYB/HO3
rQYhXyP3Yj1WwABFNELYafxX1tsxaxW2N82cs24/N13b7GlrNbSeqdP2s1asxkJr
Yt0dpzbR72DB8y5qyZyEj26EKlKdXct7AgcxjvlgHlXtRRHuk0OCnv5u6s1pgT8G
WozZ38Rb+vw3WGv4gzWwckN252hSf85zqifDMJCfjeWZok4chtygz6GJyMggUC2/
yq4SJ71xEzduR2NA5XZGzzYkMwkZPzZGRjLwkXA+Nxcp+daAcr1kVkOAa1YrKXS7
4z6UcAcUxYu6aZ4+oMLq0dz1DXn7BxSPLfJgUSbsqzo3JONAkjIjaVNYAaOUsXlV
uxn4AkK9fs4JWoelo/rC8vwvImZFck7tJFwpHkVRlSrszfuYmA3d5F67b+HdIJaP
5r7S2XVOoM971UNJvdwNiSCEQKKozbXI1bANINZwbB7kc6Pln0+gRIiGkf5kFjnr
oWZkZUBti37l/gvQFz862edRYET6KbQpgmCqDAxlJaI7uT/RI/v6RKLO4RODXHnR
uT4YRdJoSwdr3R1HjX4/JYaTw8yo+LRsq8dE1q+Ayr8suATUIHfMUtG1naFPlN+M
OdqiU4SX5RhfUoaKIIaV+ZRSNEjN2XJdXdNG9YQUd5/BsMr08yNg7yLrjnuRG9JT
zVIoTe3Ooxq26yyChFCcog1Vy00wlmn8ZwmSanERTyP2QMoNlXamK4rTqn+Q8TYw
fSjfDcRVmS+zYq+foeMIaANgUOcXmO6cT9zEyk7qvN9A7NRXrcpmPxGvLEyxir8X
cB3fXQDOY5jSwmf3EjPUZpj9MabYYsYXzapsSmBKOXXQzjQZ5RvM0tWn4/0HJt01
p+uqeu6UOI8jq4IJxLpv2Kvp+SX3Sn3dd/YsLkptGyzSxXMbyptRuh8lV4VcQaOS
9zXUVX+t2t99U8zyhxeqQ29XBs4OVnK+QRAHLW3SX/ht52z/GRbTXQDMiOEBOiWE
hIu3OLF4QSeRk6nV6ntIuOcwHINsSH6u89yoVgthVDqVSaAnB1uoLckfxCg1l5b5
drWDgzyzJmIb/YYZAdiPg1c1bb77heBsnwa83zxlAA/lhWHxcJl9BNAlmpi1hove
6DfWftv5urq/6Nz0VYOjQAraVj6cvaJ698dplN0MMM9p8vdiBjwKHR4aSs7aZNh5
1xF0zq5pJNk2DPxO6PjiiSKtrOLvcUwR+R72K/acafrvPZBlEfvv2FEswBbrgkUl
HTzpWdNtYNTLZ3vbPjW7OyDuHgJESqpRp/CJukre6OIITPbBCiVGm7T7M0Wjx+3E
uV5jpEThmfsVVDE0etGzvjNm23kdMZfP3BXs8IbCtKQBd6JjyawxHuyHwNiKlF33
9S0BdqEt0qTWOvKDwD4vbGjstMKvxyZtHct5Gbt+v7FYyD4uXhReLRCn4FnpO2IY
bIooO5VzwvD1Q0c0wrNmi8+hKo69mQ8fj+kCiHfRSlY8xVbmJEX/sDwCY5M6vrNx
I+f1g6WQB1yUMAFBdyQA/MiD7fhlTB6f4JMrp7VFJDrri8NYVR+VLoeLIWQRqMHL
uzG4THgBrv311R+3vB50DoRjRKVM51eTqaimX0GiUyBa9SQfEHgFhbvMOW7tQT9V
UPRpsR3q2czRDjwIP5Dehx2ImZGuaYnPB0buRtrKCgM0ODlKKwg4jT9s/4oM0Zcz
GBY+Y6KWqqzBqeak9ePwwJ+xaleXnmYWrfDejuzsi7BOcc6wzgqmc4oQlwADXtC8
kyFOM6GrTfLavuknlUN7cM0abnnqwxudUwu7Dm+ZzuYv/H8MTw6GtkmyH21J49po
A+2qkvfoKYnpc9Qyblcnu98irpNLNx3j/qzThPZeCtQL4qZqiANPZxChHwkBaEjj
zQDWenxI7bRF//8A8B7zhlxJzgzf6o1U332eaNSoC0c/A5IolETIM2Vjm7OpM8C6
af7VvHBqLXiRJnsERAVTptR1J5qk8p1zJxsnBl1fz8LHL00SvG5m4157bQxVx1uX
IHZm78CmNL/uvx2fV1uUhKMB2iEryfG9yz6g/SfiCF0x3QpbcoIKHzhS3NCI47xF
U6L6LK8hxs5PU1XhLAaC7JjG7m7kZRhWlLl89mGBaG17C48tOVP7DS114yLGvSiQ
+g4VvtYha7Ts564rmGKoBaOhHF2WXnyjpSJiWLebm62k/K1DyOQK8MJFr15D3/LN
HcbG6zo10L4NW7b7+V5Y1DkTvSoVUXOrj4S38rhV7Ecg4ySrxCmjApHzSC7W7dTB
b6NAvcC/M7O/ZkV9/dX6+2GflICngnNMEhLr1hcqSF2ANv4Nx29CtmlXVSvXKNPb
OsAOy9LWZvDP3mv+T5zFCxMmhRvIK+yQv9MBbvVvfAwvFbvhrhk2dyQXB95uSttf
+FWCOtjOUceSRAx9QeXRsKqaNKXNiRF2Tg9YPpZfIOQM95OzBqr2Ze/q3iCxzSfG
h4vrL1l+Lswan6yEUB6shNJ/ItbJFrRPz9jxCpofn2XtpqNvsHp2RDFz2ApVCWbn
08et3C8uJnLEo0IC7nFj/oDHYASifNMxuOyDMpbaRlqzcej3tfa6GdqCDJ2cYPeu
gUyEQDEICYcORPSXdItaYmN/KMnjnm440QNNV/39No9clhQ2UYNBhTb/F0vSgf+i
LxkQpqYj4TNAv69VjJw1AtHsGB1zLM2gzVJDXh69QlwsjmzgkXh/rW8eMaAk6X/Q
EpPe+7iMSUA8ZK/lhGlGoGjhLOuJsDcmjZ2/tmObgba9Qdo50M5iKTP5MeDBoatL
Bpmk3mj4TIQQ0l1FTY+qThsk0Sq7mVQwq3BsllJp0hQEMkcZ+vamVMbeS92ayyFL
sB0bA/qMl9tegJwCS77EMpuQQXbve4MkdZ/VpY6BqtzSDK6+23MLqa1KPmFe87Q+
lQEvwN3HFSd1qmE6Ak2DpgD6/150uI7Q2HvVGWUJDeffDuJ567p5QFx5K4dPFKTW
sqLZ+CGKgtfJ7jbJdxMRkeSicL9c5ln9VVADhuqXe/waS3lKGBT2/vJF2e3eP0LQ
lewPrOPwja5kfMrntE3qHNGCTQ4HPbtjnXCNTiaXk1TaWqLti63uSNLzioNeO7WN
Ynbs+5z6eU5PI/YiXWd3BVVNZssazEHoqbxKMf/kcnw0GkAWP9xFtPY8XzS/CPIh
JJ0w55Es2LT27n0xzQAmAB0cI3UDjsag5jvhgl7bG4qFDeVTsbEzwuItZlBdNBe6
5j4vp8i7LAwYaFUfY+z++ZRHoSfR5cb6KfJA0+RvSIKv/4xfMPgQZIBOkT5Ne/4v
GFkOMGN8YoMs9GYHQ72XM9vXYoONM+zu26jDolR/gOptlSdkLRHDbA7latXuCbqv
zR1FxcuYYes5rT79kybMUSXtk9yQpfbXnJuLIkq1geulSwwxBgUZSMI7NgQvved4
5r1pngCk/NmVj/YormNwsXSwhe3ALnzauTFxXgSy4I+v+EUC194EIKHkV2HzL7nH
d5TuBmEndQdE+u4o01dCyk8QvaTegC6XiOjErlYbee6aKLYxCnf2w9LNnEjKVkv4
bFNWatLmQtRhWpzHEpJCrfbZKSN5/BLgC9PhlfFpzgzspVU30vl58dfCvHqO88QF
4AEyh+Q55xh2PFByEQuyROnewJcvX5awW+f0iVzN6ex/4UC4FBQls09SioYRGrZi
SpVCEV+quqxj+SwaYRVet7yaqkCe31CeMGctwpsBeXih/4SPNZ7WkPa18P3FI8RU
iTo5ShXp3qzf0hufTdOuFfoJfAE/s7IShiXR3pSFN3x4LBSmZWNmL0g6GfLkLIzo
9wL0R3QYWlryJ8i0ga7F4S03cPNhGgORhk9kHzDBt2PXqsD775hEKIQnZDzAuOfG
lBSBqKgywa2Limw0q0LECCObUNNtVJIOeojxlfNtCr1QHNKw47Rpt4fSXNMjKQYw
vJfHA+23KpxoFk4NaFi7gDeOhcDem4IzmEcGhMz1teEqSoAUjnyaTIa7ZabB+AHo
ROaL++FmNdbuf/+tRUFv69UMxIzBPPoxGErh8y/U4vlI6C29h4XUkcJNJS24LpDY
qtrLtU7V3IjkjAwy3W+PnV2cFAa2mmBbmGJAaJxLX9bJ9vUU/dpg75TPA16YKrrT
TMlpLPfCnDoTgH9BidmzrwqWIft+Kfq3FleNJ9Ak2szwlbaNdYkay+ouvsIXoHLM
gNqWmkOUvBoqsSK1AXYC+m+36W/pX5omZ3AzDMiy86O78FEIIbfj+TyeCCVE/s6v
kSD3m3bJTgR8P8KHgAGEvzulls1IDWm6teLsPdMDewFUVyGo6r5XPyyK8KxFscGg
PmQSRxfH0rpPPd72K1E1rPNIvJSHFpf+YWfyORPRVmXRwrcchb7USgWkXfnG2+nY
6lkqfq4hNllCYRFFa/f3ENCRZ5ZJCpP2DfkXPDfoiuLF9qTCEA2geBe1gstEM6xH
T8HCfIAVxHKywo3fPDkvUSyiPS5UX+v5scSRsHCsgGXjZ0K5WLgUfrDq54fquid9
NRyrl6BRDp90b01dsF0qDcXhfuSjQSh1SLn/hFm4Bk7WaMh/vM3aw6MVUhAvsg/a
jOkMI5J6S2UwXmXz6PjrbuFWhylFcV9r17jJwo3m2kAtDYxgT/wAV13+7yudYJGW
WYhsSjPITTLahbW27lXZd0IwV+8jJltCNQwVWd32KzTTZQrjmamlc5JbG4Awjfe5
ZCO3svyl6exFWe5Abq9s9EvU0itldsvrZu9c5/3t3wf4jSKZ/KcfyeZrD45i3132
6Dm9jeSwW3zvAB4jqbVR5AYejz7RH1jHhDqC7AQzr390RUGpfvi5t0Pbc2OLfx5M
SA92xE5P7+hOFI2cfykINa8NwPlaLRpmprfU2JRWZ6HWPRadCjiLpkU2p2RVZ7cv
udDAq+O3kD1mZzebpkr3S6NGehj1qx2VWTdsYI0kvZ0syh9srW0/dmNKxcyZj5yn
6I/MsnHLLICuu3GrlFFbvh6vzjc9fr/YYbCxcOt4HRmKGhVLbsVklHi3gtgwB4Px
61y+wx58+WBc43oMM5Flepjp8aQZ8BYCEuhGVnj4KkjOTR3Y0EiiLMb15aC8v+74
dq6Kxl7/fn4lIBDnhIXyuPQvvelOHEIOlB26JEFlMXt/HITBhX7gyYFNw+xsjBXn
pfclyb1xTA8f/m1eDUXzdFiozWc2F8Rz70nKTrgOPN7DF+dDD7x4vEa8AKyq3lgo
EZWlh83fQC4wH0TPJ1iDV4jtNKDtTS8Ywllc+iwixEQ403AXjYanC4AiP3mlPE86
Uf8u737jEQbsy2doetCYjYpegwqq8GcUUiohducxYDE2Yjrm23sEIZHYhYEDS5uP
TRXrWUR7TCxE49S230vAx9jfakGFLJUHMgx5LLNpMayzaJ04HJpWM1OdBlMlizZm
d+aISrlMHAD9fjeUMfpENVikGbd+8wsebdVymeGuEWxLDOfHyBOpuMdhoyHHeeT0
hIIBjb+8apIGs8yW0tR7o44FrAISdWAhAP9C/iwmDC9qwGHlfBG3YiJxJtqG7Igs
Bs/oaKTUMMm986RRZ/pO+b8uitVbnGrzfjMoFsbOn+/o2KEP3wHPrQ91hzmPzdIz
r44Y+nl4d7DpJyWciHQFbCs3eK8Kqc9kQp4WuBT4lPbpmzoyHDwKy4LKeJPKJ9he
D+lkHMNXThaLretB8oQOjSKJJIo7KyqNsgCRD8SQVuWRdHK18pu/1vckXc8kIDD5
AS8bgAXqV8yAHhkx5vaE0oh6dxsbE5QGRl8EbS6BTcd0hOLrTzGSxX5cPxOm4UJm
i/24+oRZvqEoaxDegN5oMAFKU2absglclIJsYFpONI685Jh4wlLvCleKLE2GXlQG
DD3bNgM5vHKkLNb+wr9mN465vpHJjp0l3TfYRxpw70aIIGLX4vN+dPw9Fito1VX0
/ZAs2iIATei3Mea7966JGfVj6TPMUctVeGGheEgk+mtkVwlu9n7UW40X6TIPBOug
qJXX65M+A1CpnDtuML2VRSXFvIUWGVRmemVVfbrpv91N6VqqmavvUikM0YwnDgUv
Ss/K3C2tEXxYT0V+35PnDHDb5yFifZ9WuyfxmM5+3vw8Zc+5RHlYJ+2RiMri3XiZ
zo98/fwQBXV8vvGxqlpAddUcshEvJUfeKIVMjpcxW9cpmKmW9d36vukD3Keuj5BA
/te8no29cYX0mAyyTtvI4y/HTxLHqsgNceZjrihgTT7y27hsexqdhmqnABFQ+MNJ
aXDiXNniipf+UkGVzXIYzggqm/Wxql2hxa8ErCD5EsYHPrcHSO6zkXvO3sTt2e2S
FMKVe4OVPwgN82J1QYZs7+Rag+lCdeJaFurrd4CrvyWHvviL8/cimoOIeMXXjeEJ
dgv2brlkvlqE5F/eeCjJTn8ZOBjKn5gtQJTM5t58LV5oRxjpDagxP0JTBn5BD6Fn
T5889yHt+C/oMgbIBRdhQ7I9TA+IXjA993Dy0v0ZeWNoatArLXNBxFua/OkoGXEF
ntkkZMlfBYOXnGoFc7RcxJB0V5cg4n1qbCZQ+UvGdHhuw0fFTsbh7CZf+VqfxzRS
Mb9OxXGLPpuQNL5yq0bjDCbshuyfj4lw1ElcZAX97wynvvXI+hntuEZdES1Haj+h
VMIGbY9b2GQJ37KfqRUfFib+QFAKwEU7b6EOraT+m5Jjixm9BeuOCeVIsD8CSSB7
RRy0AbJxrt4XwQawjLxbKm/uTl8vPgmj1wIYFM6XzHKrQZqAwVbIG6OMXC2jFFyI
1S3h9jWai8gm8v7SQkGnBxKglp527Pi/5If3LUROfncbKIziWtzcQdiFOJJQmoH2
iDROQCztA/znZqHmkmuZKOUCDach1FWE3ykMzilOCxMOpsChj6FGyxGZ7sBwP/lo
jTpDiDkgdl5h6pTA25R9bKiKX21p31Y1xCbeSIchPQXFGkpAdtYSiuDuvjX/c4s8
037j1fW1E6mDYQfYAbEzQolw1ZaEOp6KAGxanKzvRz13E8HOzF/t1U/+K/5m6fa6
FC9fDP0xXu10bzSYW5/2r+2scfkoxBHdjNNs25tP3HVF4NXxcVY4g2TDZkjoMesq
GVcJkHfTMT9rW1YHi8b2557o9dse313aUy5K2kAAbCSfQgUMOBKyb010uHWNwfv5
UbiJgPmO/MWrxIJIFuKF3Y9tWyUx7K6caRrzv/j740LO8WglBWDyqfW9Rz5zO9TS
BS9BcDkMhIcl0el9adD6AL1D99/OSf5YolpSXyCsHNx33kPMkciry+wfKD7eBnKI
Q4GKltr7dxXHsmdk3dK/WdDLnGK4j6mB/xnMKhUjmSmektMS7rh/tnmpm0n2F7t0
lYRdF2bterXA3ntHDYPf5qw04w3m856n/1gW0Y+g/7yJFbfPRDHpk9TNh/avCSuw
TBnRWmb2KHC9p01HwWcpZVbUSli5D6inmYoYWxElmTPexdqQpIp2tMyTZdn3JXrG
lARgFjj8h95J6kDFJdESYM314j98jpakXQgEd8UK0MNdDkQxgLrJCd45jemrl0Q9
73KhR7/9rQ7h/tZteDCnJToOF2SAJeJDUipgFvSIJi1sl/kO9WofaqhAeSPoEOqX
tCqpN33n+bfNrTOU8cXCWOW2k9vhwFSEzUZMItRznCn3tL8s4ipkVsz/bVexkplS
DZ44pkhbJNdYsm82JjjaSDGDHQsAK2BGJBy2smuH08Iwfw6W8rBkHrUfm64GO/Lo
REPo7g9/DsWBq2qvKuNrnVZHddU5eYz8XLwvf600XVidL/gXs+04RmTDNoCuBXJq
Py1jB9iV4vDfhtX/+eTO3A==
`pragma protect end_protected
