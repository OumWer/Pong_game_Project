// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:01 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pEm+2CzRNn4lyIGq8GtkJAW+oyjn2gyoSgZ5JfXEn4NvlD6KK7MSFtIEBS2dtp4a
bxl/tdiO7bV5NJhMdV86xxNn8ler/qDpcsChUrTmvFbsgNCpc1hk0qGpR++W9mQ8
l5bpCgTAT5l1+2BwRVjyVz1ntaTXy0W+qbzzKVK8N5Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12960)
Ikcj5P66ZHNBT6REywJN/jV3OQFJtIXVJ99KkznDSVDd7X+joISEp9b3s7PzvBnI
oQ7dzxebL7pvMKwQcHivDFHGsJypA8qe7c7Gf4r0+4nXLJJGUGTAY+yPwc3awGaD
qcWNIECU6W1ioL04bJHvQktH96MyrYHbILbGQWoNMvefMg2PVmD0XdpqFGFTEove
g+Cn9+Y8BaZJYxRimq1iEEGtNdVzTws0qNhhpjQANpCzcxElFZz1I4KCPV74r8/G
9jxQtYnkB8THfRUYWGynXZFxqE4X1rG9eneSZuBiGdXiDaqwN6T3yijKfBNJoVZ1
unx+dAoCYjWzXL+iby39UnSdqJSNFPBddEH89ceOVQbRswPkNg4kuKXfjjPhtA4e
H5rAnIFtmjzifRKEN4NjT1O9MOMJfl1ye99ocSdzM6NJ6IvOm4EnxhZZhzve6duq
ekTlEmAdkgB7s9AL4tNhlQ7YdKksSKCXwKXG2aXKrWpLI85EWL9tFfYM78ESVqFH
Wdi7xDpUlSBh4n+IlGcihbac/J3I1h+xMv5hU7DFveYm8A2e3uWT0lxdo9tSBcIn
mt+NCFgAVYvnVbRxVyUjL/uTCXdyqupctBfgxGv0n0ndBse0libD8498uHj3syP7
8j2AVbHcYDrmg0cNiGkjRdiT2XC2MlfHkZLRmm5Nokv/fvW6l1UbkqTT5UdqyxoC
6O+7YYsZxYpo6lwxiqQWgSrVhrKCrcKO1tEYLbJ8jdJoVJVkB53dqjN3Hdtm+ZO3
qQ3trlpd6eAu1GtZaQ9BEKSEv6lET6JWKK/ScLitv3EWaQFF3gZV2lrHavNutxqZ
fP1pNKoyOe+JQx8ghb5CvtW9UOKZuAqRvQdqaqtut9+NZAjerif43NfgQ5zhegav
Yi03LxYbkryjqAontE+2TaDnmiDoOF5imbeYMf68VVUb4QJxb70xQkHYcnADi0DD
/K4GZSs58R9NDydf0UFeZFhMtAFrH2YDJ9XL/tlcncXw2MAWkM26n+mJmkSTOjXH
3e72x/3hT5QuEFuWPaUwcNtN00kUspjC8TKQTXmbKuZTCC4j78mEkX49sxUDclhY
LL315mCt2InrLLAjmVVhJsq+6ja8cTEuUwR2jkdlxnLYkACA824r8dKQbEYBd3MI
gcWc/vBdg2+uXwKlS8i7KPfPgVe9msjqO3ErDWIq8Fioytqa1r6h3Vmgjo5UOAM4
ucFmCuu6IDdehueamvdLxWx7hVZdMxROh65IDJ5QTTeOuv4etLsYAAc1RmXApoUl
LZ42vidTyLOUP2OZ8dtw/0PPEzDtUf/6e/l51NRS/D4K/nDIYGycKiw4NBJk/G83
UzSXFcQlm9jdptC1HeQe1FwYUDGS1zOHEJ/kkp0q7JZCnTGi8XJ0Nh/gl7z2ONiE
hUC9+ojdGnx7gTUG+YZgsc4QDMEV9ku5W7EcV6f8vlpX2RszGGRaSWt3cvV375nv
YwyCBWimn14+33lIxOCkdgYb59slRxWRJH1+9tIhnqULpKqJHg0lCgXOHEY6/vjP
V96SurNpr70UldcN+haHNVcrVKIhB2PPnETVuvRIZGH2bjht7eWF2qrwQAKA1rFC
0j2lNF6vPunMdbzifR7J+wqqdDi9fU+njjNa5flgS/AsLM9ZxiI8IF6l36gZrrCt
D4v2o6GuN/RnB/UeMy4WC7BmZKLP7GM2YLKnB6ao7JpKDQNDCnzqI8FP+/9ZmSMB
ZQ3fhz15wqbD0GapMv0Wm1HA3E/mB9JfEHYNlPnS5e/bA7lmxofEcmBD/C4yaWKY
GSBXmWkUkYKWjRyNnuzBb1UeLj6GhJZRBWM2efQpewaGxEFFD9n0xwWHW6KwCJ9P
9M9o0n0SVo2NlrmtskxazJ5wZp/MuF8Z/YbXiPYra9iy02y9Iuos2G3cEvXTRnwH
9CpwOEORVlfeasndJ31gH9Fy+35A5Lsgg5c2OGmOcgCAImnm/m3FMiVCHwNy0Gzh
Gq58yZZxpEP3ITNGa73noWEorJG/zdbyLHa7iJSrTQCrNl23xkt91q2Ntw1tjpf1
YL2w6Pa633ZMVlOZWr/sn+xjqq0kvm6pgoc2KedBtTakMXamo+7fSqOjPOuJoK7j
g59m1TTT/rz1qib2Hu3rMoVI2L/OKrH0RuA0CoQJUdj8D0LBCWpLMMeFmxhBye6m
MoNm8XIG6ZLTyZwQuLlbt7M4xkXr8osm/gbIXJ/bgFtLsjrCf6TB7owDayVYMWHE
AkD0pVz+JIz4GYrxJaZWfx4VNQkFjlyQ9m0m9EqGFglMIFzPFHSZ4x6CB5BbSFqh
RVElf2Vm5WAPde2oTYS/uv1jADG263GDF7R2lOrBaiIxGf8X5cA1cnKKnFEsNolt
SeAOE4JmTiXQkcYFJjF4jzau9+8yOmBojD6uQb+n9c1eWgtWAWKPWTn45SIMqxXv
37xjZrQQHTqV0rJdVDpQipHlf68JppXlSUN37mLMPhTXNKF1MkCHUceCxkSD0+vI
wlhO4q3/VrBKqcOOJ6ZSrjQ/j+bCsRxa+HXnJQvN1cb7Vj9ArFu25yf7GZ1bi1bo
g0WHQquMOMShKwaCsEqiwFZXQMUfSdK6HYJ28C5L/7YprkG71MM/XZEKGCcJqvU6
iJJasUABHd1T5ymKKE50RQUR2drcXZfuVpi/LiI6RsqBEa9o3M7HQZGRLDjTN5s/
43nbmNyPpZ4kmIApn4rgcXN6BdHFa52OnmIHx6IxPDnLQSSldlzuC/o+eYPM4hhE
LY5K9f1gY8uftLxUrbDiQ9LjBi+6ZNuBOko+zr6bNfyUZJVTiNTBV1xvCM5O9XCt
PJXEmvqH92hmSIlr3RBV0nWEKVAG7gRPzDpuUeKV75aH3kayLgUtXW4Ldty4kk7f
ZnqqvMTs/JbTUgiGZ34aXMtgTuKV0i0beYyRAxOywWhjh82bgQ4TUtYXDjMK/8OH
1C821UGD7AKtlpnMiP7rY6gkdqlHOLQG0eZEnvgpg0FjaW6jkG7N6Vu4bk46L/NE
rY9zl3/NPCFaNE9C2fiNR4JBbCO+/qqacJ9LaZOi6Q28gFjx+BzIijEci5fPCjBo
1vMjxMM4iGoOtkQTzKqTr10CWc01Zd/g4hF7QTe2lW72A+UnyNHK/Run0KFgyIdi
UUHSWSKV6EhSoK3JqhKWpwaMAFkoZr/sk3qWiUXKzleG1OfLDLVV08IOiAKQl+CG
DZCC0TN532KzVxEc53+jhoTAve2SVusyb+k8fcskVUY2drtoeIxAajB0MNtb7z0w
GHdVd84zCqCFI9w1pMQ9YieE+BjK4H33hjU5U019IVYt/uGy3g1lYombIQ5jl8hS
WsfJCk1BCcxghKYudPdBsyZKd22qpY7UKthoJRKd6gvj65irr51f1grg7PtnjUIY
nFrXdfvQsXHD1TE8WfbIovqpqEF7M4xMmP3e2JF5j+z3GnrH+Qpc/K54/pFV/6b0
7l6mzv8zznpL+Rs4noeqWNtSVa6ztQt92jVBs0BubiqNCJT4GxeW7Kmn+Ampmwxs
JD7o1zS0V5TU6gLxiT28BZJln7sEnZp0Rsh1Q109zEvlUMoLGdbwZKYV7OtPTFez
OtuU5Yo+Xbu8Yl9/fBbgDh0VUGBROSP6IOllE8gBc0JDX3L9ajxdVR+gF7GCkGSf
ZQubufPgAR5pQYXlcZ/hFAv4XaZDo0/tR4llMQgWnp+DA5S43vwUPWaMiNJCHI5o
TRGsx0xhHoIcoiK5vvVUuVgtxoMXKT+CNuQPjRP1lTxUy8WeCI3UThqLIr8QcMgA
GnURD/fVJ/zZhOxacseYZEyvRyuzQfzjjHzc5ZfCeHgta+Nz5Uqtwr2WcRRozGw7
oFYc9gkw3WK79e0GcTi1Sh5BEnhQgORvo/6NvIC2z2gOShCP/5EtZkFi1lpkJoIN
MG5tw3ipypaGIxQni1STgbANUK0kY56k4J2rja8lTGjlyMbgoTBJJ7bQQN2Iiirl
joOfuVhDL3HMwmmSpit2+E42TeczJm565ZznaihDN3dECoGbXcFZtdbZjqI4AeSw
gUZwFTww3KD1xWfJricm5VzxCYwpp/7vyF5k/B//Gm4DDeNRVah+KgXtFZfqUwdP
O4PuqCzLIxD2e7k2EQub04sz6CaoEaZYtRd2q0tcsp6MDKy5mdUzoRVjRni/fZmr
bYGxeFX7N5g2jgCTk7FDJTNd50DM0an5XWm7b20hHq9heKccihGehlZf4Mh7iB4/
tD9ryGHk/VOq/0b3fgpjd5qcSUKhf7wVI9hmelAG2/B+c+nx48jK6Km5Z9TVZO/n
MRN5MnZCpAuGNT1pNfH9ErQq6Y7aVx5A4So72ZilrigqXgoeNhAU8881+as/eyRO
R059/PVVtgME9UmUL4Q7asZk4BeL0yH6GU0NDNK452gf4f1llBQ1r3HNhUDZl0zN
Fb/o4549hVUdbjwKIoiyC8IpFOivziKPuX6CXy0lV0g6oVGx7QIhjPaTH5pR4HoG
sgQWlprihlkYErMV1DYZCHSSSHAXjOPCdc6yzFulLqVY+1clhFHDO4S5C8S2IIAN
tALGSXOja9LU4heOKVWz6bCzDuLOj67tx4U7xVVL+ZT3uze9EAlt6zyDP8L/JcuL
IE3f8/yzr0FEJvfs1a6iDU+mXtSoyAND3KNHHOXjigyVAKpcVfkCz+mHWYmx/heL
ZQm88JY2zXUW/QZBeBXlf0i+UWxyR9BesBVnN1/LVGzFlJ7lrI3kRIFDSIltwLn1
0r0S5lYWgpif6IFqEzdTGtWvekEmAZ+wX/XJUFILPam/CAqDgQ/fZMIIO+pUoN/R
BA3q+VKHAMcesgyqEbbezQqw9Uy7TqcXqOYKGJ79QCvYgO9uHSyqfg8qhGGDi9Mb
cGCv/kDtv16Y2gi/c0IUng9wh0+ixlEH+7/vt2pG/XPMd0hcF2cparX5SVqWqeZ2
cO2IkEBoKUuoFN4SvaSk/MXl4crts6Y4PlLUnpVoO9xY7qcugS+GRu5BuKSJ4iVf
iZ0OCuWQEaQkAWXjgIF65AYRlvx4vLHP49/SFPi1tOb6o3T8QplFrcPLUOYX9igm
F+nqH+hT6Z/XlTh6k/cspKp3k9UBh6UkvJMHNH9cHPHvTWXH9H5+0qtxDaZ9ypQc
7nWX8UyUKQzUtbnixrQmZ1eMAWnteRP4Whz4VUdwcXQVNyK3SXjcB68S+VHWVEYQ
kldDoPUbDfBNFWrItuuSbQrRPmhHkP9Xi1YR3gOLNHqQ1AflptI7OYuZlRqmzE7K
Pl92h9j0rK2+tW0OaX1Cd6KmE5IXIblYttu/gsAS92YoAxxu7L6LNbMCFKhAjpbS
X0SWkWMmzN6oKPs1LfO/iMuVcI3v2OdsNqcnMWwBmH348k2xp5xxFB3pOcikQh0b
/EXZ8//d2ruFMpxy/gaewdjkKKXro2PDkMY5opGHJAl1S4mmobtE0KCUJGcZ4meE
hl6OqMDNtcZZxBMGTxVDeMi5O5QhXDQ6MlROo5vzHxrkE/AfxBEZbKEORTAOk7Hu
piJf46wJE/N14BYrueJdNSIH555IZhCBnnT9pBzk9tEAifWoK5+nzUNujUN+6oaj
389wb+DbIa2FVt2ZSEnnJMJ8cz2tDALHJ4zvPKrpwUNA9MFgyCNzUbCKYpNcfZlZ
OuEeTHyi/Tc9a9ggCMB3oNBrtWc01IA/b1SS3JpsYr/AZU4Edvv3hmehjT6bq69f
0zmRjRCg2pwGCIxMzwR79zhbU5tmktYN1ffsQybUjnEnhHt06/84IKkkY2FiqBRE
gt/DSjtTJLoVdjxl0+LssNIWAe9re77aTmZCF6Jq767oYkZmBJu61r48VXvyKULt
BH8UqEI17jH3+j1Cpp+Cp919viI3icFvSDjoCaIuI0iUNe69CSL+7pQvE1OFHFiJ
9CZT2aFb3Y7AD5Vsxd7TCfSaH130pFZWSwZjcgONEoexyjUMX3h7F+PISalr/pZS
io8dP4cSHOmZf86Mbb/+0SxFaZ1GxEuwUu8l7pZtDjjnK3dBRMz9Ezd29C0PSat1
WpzAyR+ZdKVTk7o0WC/ApbTciOoJud9mnIV/TwgqGP1IcxipJAfldz2ckzl9B8nN
9QQE3g/qOlLHgGTnqx6oVA+yNCActFhyoV+Yagbm66yvTEaRVnwlfry4H2dD60yV
LQ8EWquA6itj66hMTPxKaz9IFoQTJ3Cy6z73Y5toBzUJovbiU4nfpcpxdhvIg8Q5
JQawfQXBr2M6SU6QlVQbjr5G4ppTb03i7+DJXw5B291rw9Mp+6gHw5eXJLtVqcz1
ila3zArZzYwKKsXpC59BxmGgiVQfHGU2PXEWvlFSsPXi04LXOBX/NrBG8lyVTT4H
KoZM+M8hK9L6jEyDi+uoPPcthjgCAVcdkNOAyQxdxy6dgzCVA38oqP55IMsd9W63
fbUGgsK/GPRbgv76Sk0PdCHNMwJxhDfNYfjUfAd6vEcRlgNLGgs7J3zj+yf6jF6J
0SlzW8nx6gwt5xm0F3yXJw55SIhYeM4zjoS5L4C1hQl14zM9ULn2NOhcfrUD4aMD
JEkzb4NvLfEHv3ZG2xgnkHYnWo4jCHgRtEZkvysxr4slQTgH4YBJwrYxtc7e9x3C
FIw4NurB/axKo9E839qezQH8aEdxmvpsI4O7BToUe48yChUzS0rNH/CD3oURlayN
Yt/oLRObnlSN1kReImjqZ6fgQQTyUA8R137s0aYj1aDPkFwbeEHWMryvoBJeEZgW
wPBCr8GccYlxQa4QSjeDjU6rExhW4/1sd5rbmZJYt2nHAM1euZKWlctSRAijpe3C
YIALehKCzA87oS1vecz7QFwsv7/S5jie/Y8qFQ6m8s0mqB2kUE/wIpXqXHUpMR0j
+MR115s8Votm0CytSMayLisslWjWNQuo+W+6pQGQhflYGwgHODrM7QLVJR07IqTs
3zV/qcx0BDGGkjFXZsyZjDDkfFDrLosj4uGy1Hoxo0YU/bop3xLu8wzpBTRa0VLK
4qLGnvpuFWKrliVzCEolnIcZo4+VsRWhf4uSPT2LRnV0Lz7Y0Ca7Wxf/3mSKJcn+
yrE+aW53Pa/3y/tPai4Rh0ifPKPPgaGxFaFdyCKUCbZ/QE3RWn/k13ybiIpFgpo0
YlxYAthTkCKUN6//0AdHp7eJB2+1Z9GXVBojzDWtZMtOHvAWw1U6wl8pdAdV//OD
v5spQImD0padCE7LuM+opCcLNM2TKoxRhe7sifAm2nM19POWGk7gSic1IDPGh7P3
EbQA0ugzNd1HFINP/ciJ2+M6/E49a4idgc4YVT09Ff1otkWD3sqk6p2u59XF9Dge
yh3gCXnivoAMTt/m68m8SplhJzoMtA8z5FkKnv32N92rdHEnYoB/aEornQN73FgO
rTuoKWhLcR+09vIbPPIeRxzNjKyPk8Hlc+6UHZpA1S/jltWdIDaBXC2v2MM0MIOK
2X7vUol/90qLkxA7iKkEHyEJfrWe1JepM7BnSKngdSucHzMbMJXXeIQWaG61e3iB
YILcvaKoUrtLTO103K0b1BKeGtBykyqLk/+W2mfm7wKdlY930JM9I8bCcmv78ZRn
tOKIxCQQ+7/T8rvTlu5BQVFkniJrcDPqLP4dAsSIMdy9rrpVs/qR7cOBSJLVIZLX
gEl83CPhq8opKv79hGRg7DrnS937hNXIhJFu7d0XeFyN6bVNXoWUz6h2shue5+e0
/gVZDqnNSsOovWm9iK1XFihFDRyqq8qmIn6fFGwp/hbC7x4rSI7MUlm+uUAO7/xo
2AM7ccUrGb5owsLAQ7RwbN4TjS146iciQMqKSo+NREvDrje5j9WPo3wIVoyeAv/0
rZp8hRr39lT3C6QPb9axHX7BlpmPQdIpHKzUzXAIiyw0nknAIvJDbEgLSu8uiMOA
Tl1PwQvmP2fCYKBoRTwgt2TdGEQscltLzAZH9NY8GJpqmczdOPxRQHNz8+yEp8l9
ZrwiafdB4g5DLCyJbo9Jh5rEZufwOgAwn2DPpyRVf0KyAft3HGFdSkU1dp1M/uVR
dEsfIDOKznDU95yUCFzX6c+vo+HVgzgxbSkTSMYzygRxXbNsaWNkVAzXr0H5quVV
pgYxpGJG1k1ycoSHm3xau/jpU3LF+IMODYpaO4NQjTpgdapT+Ie+/HlGN9FhYAd1
hGRNJsLLHrLSq5p+wXBfZD2Jz090VV30RsCc5+kxQxiJZr5NtEAI8Vz8igsRsck1
/QEjlxgeSRgGEsLt0f730nSnmCrS1xNwiphoLGmjuy0creXELwm9XL7OQK2UNza0
7viZP1AYauDyZzJZ3146u6WM3E2qgRsmD1l9A2ZX/mXAxRpuDknovlIeJOMtDqNg
2IydehqpJ7ycGohM5A0oKRMQoIeB+O78CusmGX6+ORUEQP2tk4MkFqKI3MWyTVXj
7wjmD2nA6bJC9r7jhU/q5+MVGyOnU97ZK2wVgz+1gHmuDr5+s0eu5FUH/UCEgqta
ZrsWeF+ucUdEEovT00ot4KW4+Arqty6/IUw+4EfO0BJvWdggzDt2Zy0GwP0webto
BcA6PQDdAdQHEu7eMB7z0gzSrfXRjTeoyO/9rVDJ5j9YXz3Of+KvnpTPsH46ewTK
qK87rdrk9Fc4fU+F2wdmSSAqyGl8A/BWr4htauz7qKszcd6lXzMN/zwU0WDyUORv
Lo2huroNoKD1v2oLSg3kediV5ZsLgY/HHSe40zB6Jlb2HA1pDem4RYA9kGMwc8vO
6Q3FV8RWb8MlFSU+TwOIXkKLlbBjtCjrWNgLvr4Y0cKvHuEiEx+r2m6VeD5cSAqq
Wa4PIxp6J0pPjrnaiv0NqCmwHpQAWP3uradEElba67pePm6RzQq4iSbaCXVJm6sg
9vXADVR80dQ9JUOIjTYM4mGrzZLAkXN6NeRXEnrg035xe7vJkgI96lynd6Bezk1y
PoyC+mjmK8rWWVZPCPmFCIOjXc96ItFt5mkCw3zg466/QAgLVDyYKy9pn4vKwfpo
YaFrDgb33Wkeld+tersvYyUena7C/AXpfG03K8e29C3Bk8PAtAdGbs1eqnIc4BAu
5AF/H9E1x6Dx2tGyUQMNWJKLthzWvdMM6Zmeu42yZElSx6KFnirh26SL44KYLzfG
sbBDV2245ca1K04rNZUm0DVw1ObnoqmXRlt/chq4MS+UzXXFoyaINy+uur5bIk7X
JQnEc28om5sd1Mby8OCWuk/snvunI+ACmvpA2T04vTcPXvs4rdkjncFUiJ5sgBCi
hWc6esUyh0f2EeOPy55yiEVXoe3VKErcgwpF89o+DNHfSU7lrNvdYsXLg39oo1/3
ZFP3gJhQpc4osGt3Oibq61r+qY6pXH3IUwQLPr/a3FeEfTy4CamLVRJpOtp/oo0S
PG7Vlo4e7j0M9Us3sAVpKpxf6R0ydK5KNwbPhyKZrvGwPPXgl/02F6sMdAhB8Pkl
JWS3HNIPktf/Dn1Q21Ou6JEN9TAXw/OZbJoAeCgV2+gYwhlSEjR8G7mG6qkem2dM
pg2R1+vnjEPA3ZQCMvn9DB5z//COC6Pq/9VivfLgSbkH/dbk6Gi1MoycddYLSAJK
+NpmJPHRIUfIdhhzMnC8koS2RO9lq9N2vgpwLGXGztz5Qtsem8bWqX3F1VBb9ZH3
Nl9mBnMoC/4YkCOsolM/Yc8ZR6VQRHOcofq4E1bExtSVzcUbfxRHK1I6fYBMUW4f
EAiZGqaKN7KSQVrp92GaDi3lW5ey74+yemJhW0x7+ze1sPqCPm8ZqeVuhBo4WG0j
oE1WLq4uAmSVw14dFbTZxj1dJ9AwdIrhWCx9Nq4KZ+lVY94yJV8fpz2mvCqgxukN
f0GRheggVBL7n84pPPtAfJzU7vthNkzouAtQyaODlL5Y4eLQNkJZkPCSwT/76cd2
P4H8mjjU0tSUYxvcGCZ+qlXiUDdXkX8D+ccxSJSYQszWCxY7gl6utytBhBbOkaMQ
FGCGLCAXw89BUJassJjjZEIoeACozkhGW7rTTRJk/f09JOrvdlZ1wh38aIYbKWct
vPQ5Xq9rHigH/0vJgL/DGlO9qTXD+OK2Pr15ilZnhsR7LDQIuhlu0anNX7UvNcxq
LI5y8/5GBVa1BLl+WN11Qm1lqEZ7ZZQxdO7GqEKHR5ddwZsf7bDIARLUBobYF4Xu
8zt9lz34Fiy62tv6cK/n3JpRK1ja0+Z+fhjsI5SyJeNOtDw4y5P9hFeLLs0g8JfU
STSVxOEQ1vm5A0W6rtVU6SJQM7GHIzfITDV+AXXSdGoR6Y6ixQ1XjH/RldeIyy0i
XKIuQZyU5KAphoAo9DvRhgozwxZYCM77xT+27QeLYEnqiZ7llQGKtw1MhzHXg73R
5RpCaYLhBCd98dxB4gJ215BYwE3tqYtzhPLz8lGQ06NuIccAKg99lusuvvh8Sc1K
SdhtptniClfTU4Ix0O8tsxANaNyrOsefJzDsx2KVcwIkJFG8wkyehau40HugDcEc
fgG1xAA2l7adQ9SX878ZPLPHOMRXYKeakG4l8q9esjykb0zL8pIqNJH9LluGf1X3
aXbReBhMzqyWx8z0WqjZ+N2mCwncrUZ9ZPc2RSUCcINIqw99d6TPeOsGHre7UAOx
qhn5QYwZR0NV/GMUVwBoLCn5uglweafqiif+soCsUyy67zUGPqsyk7i6ut36E62J
tUIwaTHLm+mDgho/VD5AwRkcaLokbxHgxohuQWA0mzzfKR9+j53uo04Vmi65lG9W
zswirj3eEnl0wF0LjD/SA5MFfD4OLqV5s7agXxubKNmpW6+2yh/IPaWC8aoK3Pey
01V128Lh5bA4E8gHJMNqjBZLr5HdRzioy9g9091Tyz8tLsso1OXNC6WlY14bec92
T8yN/VpWMaYk1LOFCHeB0DQWQp5sUHMQ3k2m5+C4f/fgjFCPmB5ZkdaqaLpkkhkV
eZRN4D5Tb+HTlXX2cnKu6CXSf2LHkU3AJMei5TOPptimUim/L8lasBWqSRflOt2l
aopNVyxqxZpx93XpB/DdVnpYojCgu+ymhIkdVcHhkLgNsu91lIBKRTOz2AG9JPvJ
qRZq4s6PgkPnikGclgMsQnFs9YqfD/ykRnbwDqr5djvgXC/egIShRk1+uf1UqTCj
dMQSrS3iTs0SymErX0wXy5VWYdpNCWepD//8TZh126OiDEQATEEnVDLEiyjl+V/X
cS2wyPppYrzR58fsZ+uWdDNTzwFaHlEPPT7+yBnngSLIcuQVjQV2KYBJ8D9vg0UU
GCukSDp9FyS/TDKNohMofvcHpxrQEIsfDCA8hx+I/nyd/boAujRAxlwdmpRkEp6W
l9LDj/xzEU5UPRQ1dmzuL15n31nw6XsLmq8Hb9GAMpt3NeqviuxKMiRcMGo+sJfS
kYodTsQP7skLbyNbrbc5iBgEdMcCw1F8mA2IEy6GHRbBdGQHP5GEBw6ZBUtRLwji
s3lMGhbQWsZr0FtymwIxSR6T78ypqnMUwMLbrkPvNNbmFKmWrKXOVyLVaBn7BOfq
bf2br6PKh+HbPy1Rd8YyMvkPPG44ZPy/GqLpRHX3czy2+AsbOhpw/azYTvR4h6fk
4oROl7pW2uh2uRb77SsWf5I8sazs+kKXNsreMD+XbOFdYS9fRuzGbRBF9ne5eG7n
wSmRGuhwu6A0Y0i2684JlSKgDfQdK4sInfr3iSx9DLS8jwjgvEsHg3/0rqCd30wF
R/Hi0TWlPpzy/PkZvZPjlmN6siNZV2L25FaskJltv/S9UKrpznmRJjBTRwH7K4fn
NRL+n1Ww0DXI/Ki+ceXJjt6dz8jo0N6F4Cu+s0g/BKJFoHCyxr2FkaT9RCqvi3h3
cu6TpO9PbzY8/mU1Su/BvSvG4nNGUrW72v09eRyaFvuyDkoOPUHVQbirMlGZ9z0y
9SrDqWcrcWXvQaXWrcapCI4zgm74KhIHWXYb0C3JQsqYOrMAMTBfZ/UJH+L5XtXs
l7zP5n6NmnrcCdBHXbDfKAxpsQt6rPsHvdeEiEnpoIQRmhxEcFPxakl3XFWCT6rt
ydhgfiSZfg1QAwFGEe1MnhS3qxrAiP1xK5xsel41mUoQTqOXF6eVRbe8+taN6iSN
J3i+GQ14G36gLHjENhTYjtEeJB6ciAwAprtL33bUgOI9TRy7CM0edKuuq/G+tiim
s2I1cvF2J4JDIK1nM4WYoQ9O0AEcXO8NmzQXcTEgHs3A56v8VPR2l+ME5Tp10BLD
6bYBRtWXxq/NZ6Dtic5HKBRZAsXvQrP/7q1qzwMDNrknTfgoRsKIlDgte5X4AjEe
izf8iJIGzT8UvcpCw4NgSgwLcNaI2Pf3wOy4XK8Uk17vBT1Qg16ccHBB0jxXaLwh
Q4PE1Xczp4rCBrYkW6VlIvHzeWJzkC7AV8+7ANxuwhydrgtQDSXJ25iAc7L72uW5
PE3MB2D4FgBrUbFXmOTuiSpkbQVIKHkX1g8zdM3KTJjgSYa7TwMRjdmvLgYtbrcI
4Db7aHUWoNTg2iyN2FBDFD5lXpumWnR00KgzxKec8yH0A/b2n9Js3SX/9q7p7Vfc
3hDKIzIlvwX359IyBbTjFGoU2E07HqKmb/R4jKPoIXhVP0x6sIm6+eAGb5LknWSl
rT1NdkV7rmBw3FOF4qRllPUBMsNUERZ72jTWu3sfRQVRL3CEltq/CpzUhqhl9wV9
CUln6vD+vdw7BjJTiYCF/eC/akh3NmoZDOQ1KfyH3k+5Ccb7gljJLu0PbZrSbUJN
tHPucWNou6xk5dWdFTPCPgvsMwzO54xWB25BeseCGfwQcNWxWf62yk1c0eT/GCXZ
Xh/1daE1CA9E2KjxvHRlUv0Aks8akTZVJW1z7gkgRRsmUrwJgkzzoTJMlxXU+kYN
Xt4WrfTDLza+g9X6CFKzwh5AJjQTirwQZQ50tdI3O7n3ia+duaYO9SoGUuhIxvHO
EmB/0A5BDUSiPTTlyS2pv2ad7vsthHjQOl2Yf2zjconkGaPf6lMyNAoTsMACs3wn
W9XYCe+LmwptzOaOikP/WIy/NQUzNHU17QLrKujGF9l3uweW1dWXwKmV6PwlnRz5
xo4COIc7sums8RASvfrJS7TmvJ51CP+uy1EWZbKDz3rEEfsT6B0BmQJ+BA5L/uNZ
JGs8BS0kl/16PQ6dQ1RVhZQ32zaqhfwrNczJ11q0jwu9R3pbXfPJjjTsXcfWZHTD
1DM3OrKhtWcH6nPw/d/zCQjqgtSSxg7ngzckFp33mQoQ7K1XLXsWUwRpQ9xBpTlO
/DgkuWr/hMZ0MiH0ECxzMmBOUjvJ0YmwH4iXtiTtonjHNYth0nZrQcf+nLDSg9Jf
RUB4cngBOtvpTUtuYQIGA3d9oYrJXr9yNzu/JI0j3lKJhTcJnn+TWW945ikYbhw5
Sf49FEPH2ceq79ynXyyCUIVWPR5yRHfzyMciJhBV5MW3ihKzsi8UAfSQQW3ZX1Wi
SSvdKUeorhTNK/O2fL1QWMrCr+3lptbSsAGHx8KLIZ/WzSHnBxbtktDUGuNta+vr
93PIZiIVzJpxpViiYd/X2RW/UcVjUzzfoVE/iHkNYahR+JDQ6SwTcYBufTj0c2Ju
J1ytCilD4LHION0tDDmB7B4sTgC7m9G5/Xb7wQ9y0Eh4gKuDIGWiMCOFqinwAtbc
Hk6zPIemAEFh2JVvFijlj3/47X0d5wzUgUrmC0XTDlHE77cjPxpRV4b2h24HAfsU
MQNdWTmohMcIO89ripiBxseZb7H0HTTX7WRcFEoHZl1beMnKjr6ytHN3oyw0Y99M
1O9rTlRA23dUeZRF8YROkZ0aASyA4kWm2YMkebdrLrA0qWChrj9w00N6nF6ViDK4
ABJcPOuRGNt+HlPIdivvQHCS7LTly5MaBlnRjWNex2EfsjyocJHTbf7OcPJaOXb+
7jaapINS2lUZLkpv8K+zx6CjhRXD0Fpsj6ra5am+XnYGX2+xbG1rRYYHBcdvuUnO
+QpW/l3i58/8o7iQ7coD2CPm/qhz060TeYQFLX+eimduOrEAWI1rT1PVbLctZwSA
D20Al94cKmGgSWgv/HcYqHSzZC1KIRzwr/nZFfTb/vsKYsrcfvfEyhQn3g7NlYaE
m1Si4VHkSnU1nzeajr89gT/CrwGA0Eo6ggLavsstZgYI3stP0l3ZG7NvXILLJFhp
luF8Gbo5nl3fa5pZdMXg4cm9qvyKOZsfbj7Yd/iz+jwcWb/MCEmfawfMMewvcrUw
bKfkJ7e9vyIWZynIjgoyzVrNi3+7Hbgxzb0RfhcbZWBLxVDrwluTpW+xjDQPxRPu
Spps+4LJ7fc+uJP4cIqaOldhzpShFzfO3eCtw2uZZBSVsqHiobL6kqZuwQB1AbgC
MlyuQoUF+ECmsYbaHUkoa06hnAthFfIPUFjQVHwyq/HTOd98M9ezYyLP9+fcylGy
dKV4Nnhxn24f98Ua7gye/JpJtoLYiQaNNJ/josJsEMUvEAGl5KN10SFx5HNaUvLw
PCG21uFYnztPzfs8AzvjY29Sb0xc4iycwxfFeymkmHBscQEOxw40zvqXwm23oTNP
gTzdXSUYkEpjrknJnZG1ofqRdZ+UNHNuTGDcTSUqtw988icnL1MCCBMk0eCBqPYO
fKGnHIIQQbjXPuThuy3mBGpP1ocrLbv3ot9C5TsVxQaez+THlWaIHyKCLbJ84L2H
mwnO5eKn6u7ngxMrlXpcEEgjm4gTvUQIKt8mBYx5t6nvJyKUM1G7RITbOdMre5FG
SUIMv0HOV3lMQwOoVcE4tPMV5hAjzTZc+zLhil8c4tQnMMrA9u5YdMOZo+vLbnSV
cXQNEWZYnbIKdrh0iG3fIVYXRPE/BDue4VUEDDF5xySflUJ1gv9Qgy7bpMLiyUqf
sZHD0s4+6z4afD9V7fHNBVH2k95uSNP3XUGNg2O9SGuEXwms4KxslMr129zrlaSu
BNtGmhUWNzKAVy+V1p7nemOfN6khOShkJV6ZFRWyF6cgyHG6it20bTgcIj51fcji
7u9t11XLm6kbv9zFGozuGxyKdv/KR5W4gPNdC9Y9K/zBjQh+onEIopYDgAJUC1QD
4xDlaw63T2QunHXQix2pMXxF5bTVEt8ETvBOz7kygdyd4TDS6Xkz3Q3nhQ18uzwz
iJHYJdyoHwX+Ek82B0BAN+70QhZfQMHS2hP6mdcwMy7ug+i6+eZB5yVZY+rR87UQ
+satkXYqODgZWhBdnsBXn8QKOPO2xPYqj1S0jYtSQerIDQtUkY9oI2qX1u6RWE4w
kLuUFzSEEz/IDrltt3Q4k4DXITegW+9JTvcVu+XCtzdErfsi6G3Vwb4rnhl352mR
KxNB2Xut6B7zpL2G3kyjlYkzfo4SJzaFa7U9DmV/siQK6L6Bf7WQ3+a6IW7nriiJ
51HVWZaOVGoj2hz5IFv0D1kVAFcYWe+MTgRt9myEQvyMNBkbTI3G3msyqFPWlDXj
YKXm+BUI3dOrbV692YI5xdFD7gIqqfa6mDJ537CrSlWKgdELVbdLIQaAtn8XJtcf
TJZp9d0TRJGAbpb9kDT+8MQADtlbQI4NRr/WMR4Y0mQKFVZuT2d0L4Am6Jg1++go
3mmSV2RfihxPOSFbJsIcxwxdRa473jY/A2LmISqOiAHXThGh7pIbCjeHNoT4U0c9
ebuIRja6o3b4AWxVOQ3viKOEIIz7JLQPz4hSNqhMGYSfrPfIAb0E86o+l1HgyIx6
soCM5YJH6B1LchcV/3tdjp5YPcohXA7I4FpTLgOKh7CqC8vi+wiKsCd1DjtSbjfM
e+XuxtqXGznpc9fNTdD2QoBiYJg4w+B2ukqcvESGNTo0gzm9yVMHqijLcyz/Yf7i
7CRnO6Zys5dt+wOVI99GmIGZ29dxk3LmFig+LC2Zv3co0u9NCC2FzYeGS2hlnsY3
GDewA1HJSG9J9u9npjWvZu7bm/nUIcSANJcVUDOSPb9S+irMuQUmo1fqTS7i6Hqh
shWQyZEXgD1y7A6qD23nSivkPD3sgDR4jTbF8JNKnxzw5yMeah16DTgz+4FgBLSM
w8A4ic9MSZ+amGicO2jBerDOVk/37N9SeDFMckv3lKnnkkuo9u44HhQHrvZhv9LY
N9T1RS3Ae1aqGft5WXQ+SziXShmIx6IiMSWXdmVXqnYiyF+4eNu3iuXkXqVL9lrt
OrTEej8kZ5dBv5mp2H74sUglET50zkuE/OdfzPxL6phKwy6ISa3L/ahvPhGEsGhz
5fQHBiK4klRd8Ur051O3gqtTEwAIeauQMLZLFqe62jiShmKrsBp+iVkHVBrabc2H
BISaYKcFIRt4jljGN2X6+tHnI1x85BnElASBOF60aKm6mVQW9BlgudkvXHnguzBc
y/CMewVJmHgbqPuNGU6mqVBkjGhmQ9I2PCfPpgCR7Gm94UVdsA447pn0Twn7dhM/
Xg3HAxuaBm7vx5H21QoLywOGIIO6ksHeGjj4Rdng0adndf9EtAspsNHJUYc2SLEP
B8wCDc+SDNIT4jLDzjZcXqXjwTUUUNi5PtEGv7yt4/SCdtUPradjcbK2sgnt4X1T
BCdlt7k8CEy8jyNQiw+PfGwYBdTeec0H8OXVK14WZHFT1/0jWSoQzp08jNMB34BO
H2138pJKmFEPP4x1/IP8lp3RhEKOizPIslxEqGScgMdUPPrkqHcJAr3SRZSIz3U6
pKO+uZVFoIHl7yZtOc9b4XkAg7PbcJ9VNXSXj1UtALqe/46vVTTDF2dkmwRw8x6i
Hpkpv0MZds711mJHDWrXV6oSxN13GzlLfrODNWEtYtJv45ADlpLIDxkqSzvpKL2m
YSd3s8V+NpZ0psEqZs7AnvRZeTdZWKdXZ49bIIyhL77HfKxU5vgZBe+pedvg47C4
d6ndT0NrYMziF+B2HPeorK+mNoJaS0zW3UCzIH4vOyMOaQR56AAxr3XSvj916PA5
URju6PfDHolk0jqDA90aFiMtZEOmqt7aGtI3E9iMWzr3GYW0gZ3BJX66kmEDh1Rf
pBuKT1D70UPLmhWBCpNdSKiQfYhIs6TgjdtdVI6s8qszBuOEoDdWrAWroRezxCln
JwlJ+MRf+Yoq04eg6gQ48LmR3cqbdzzswCQoMPhWXqTKJNwQtrUlTkn7gIQkL/SC
9x42d1qZ20WiWCekfE3M0DGB6stZbulvTbCYlM9wQ7IgaSnb3jpx16f47JgAw+5s
h/ytFc3F+1IErjO0u8Z+88eBN16U0yuy71oqISN1ufZV54KmZ3wBoTtJN9deahQC
DdEYz7EodfK+CzrMruG1JIYnDdNLCNNj0AHrSRSyMG1Z1S30yPeEyrWy4NNG1mQu
5A270ENdQxaTJVhT9PJar+PMG9zAyydmdCMFsUF+EWnsvQjBOxdb1G1mm2xbABtG
`pragma protect end_protected
