// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:01 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Vsdm67TuWiSpGQ+r3LzpJDwDQ6BicPoHLFEVDBizbddmEy/iKYp/7jt52bNss2Yp
Vqb3cQMDXHZQIBkHd5l1ZQKzka2G22lxn+jTl9VJZ9x4uKOVC8S01o9SRoFlAz4A
4Wr5LEuJSGM6zGLfxBSDlzdC9QuajSEt4bkGym2IMSY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17728)
5Jkpt+h2U3OckRRJ6mPw0jd9ZUwY5qeHyXOrFQ52gxqbZU6vjrx3AfvJCIIV6A2R
Xy1Mua9f73lqb3C1t76X27UbqlPKL0ve5GUQN8/IdoNaoENwwBXV+dnZwwchW1+7
pTi1wpQRGXsyt/ZiqbPF86kQrFVZEz874auUODgizfvBdzoQ1svC0YZgslHXVUTc
MGM0QX9ChJlx+sEWvuHzstPFZWHZ7B8gALUWDgzAKJauX9a+3PgSUo5T+9yYYbWr
yUwAtZTGU18NdPvOxmlk59rrnrV41oC0dh7N4Am7hVGj9b7uP7j9L6REa4mKwLTo
fjSVJf12O/rv3NZrbntslkvp9mvozVoRlUg0xXBXndhjqRPG043r3bsTiLyLytM5
dRJhiZ9wjFYZ1pNTjl6kj719blOKkiwKTYF7e5AdC27QlQDepEb7QAOyYlf0k6yM
s7wvnd8ZBjYlvsXyDa0/YC6wQL/6/P4c0ksJsGtSrv58UCAu/7wLq7gl+m7EkiTu
Um8J6rRRrj/seLb00NZsdwTujN6CAuW/LCQMQQMfG9rutTxhk6f/K8NTm3D1jPAm
U0FeZ/Jo+MYEJMh70Fz0jkaf2BCX31DxAFy5Mht6b+CdHYJSqLi3EUPPSoe0asFz
snGR45m3D22MvqNUjcGO7pKRG9u+/MELJo5BZEXShV5FLXGgAAPC4puJ2jp1fEm0
/0drPh7zGi/Jj0jffF1/9JCZrpAIYmn79yTLpqRjvqoSQWkeOLzl50VuHvlSTDbI
FbuBpwgQa9SDyCfRcc5Sg/E9Lw012zLgQrB+HciJj2Z8ptg+KyEqL4v6vUb3uQEk
7HBYCSNjjSUR5nIfY8b/1QCxw13DLlTGiNl1Zijlg/jaOgVCapEXHEhBasDyW3oj
4tHo+7nxaM0/fuKp4hwuexnv/lGUA+0xx7SMwRYRp5R1NNQ4bLD0gAVXq8YoWS0o
HsYHYAfzIQmMdH/fp5xpFBEYEwhAW8wnrCbbrOd+QEATXMf7mGlPySphzbRNEBjj
37LwIYuFJilPkhvGOWUYhCzuCZXfwO9SL9oMBrfvBllXZD8efnuyrpYgHZLTQf4D
TxLL7L3t4SrMtbajDHzerzvrOTiwxr0A63LLYFDDJ53tkLOO3QyTlGoLGYcmBi6H
ba/zYoNVdHt729mCbSFV5zNX0Ko4D486t8lk7N15KRau93LOp4gRzmrYJqZnAl8p
qA91PFAfWBMyW3OEE2slYz6oQVcEhWWQqhgFirqv5z+bNH0XHaO8O6xHeAkQi/ik
hAjGNMIwj0z6fjRJ7zbsfCcjONbReYJEpvgz32bM0iP8GFU+V34J/ThDilHbHLe1
r/kyh427bUISM2oeFRsupc1arp3QT43T8GVNWZItqLTB+5jOHYVAqRlTT5YOBARm
tvpSAb7dCpCBi+9nvuejZC9AjCJg3I4CeChitDfcWTHxOk8ECvwXk2cci3W9fnLg
uBRW9gDSd/ZqRS0otg64Wc6H1QPFgu9vK7rEYoQ6YYDds6NUGIHQUGfYhK/2AdBs
dU/M0XU6FrDBZU4DSdIKVvhTwWgcvvqpQ0PstDNJjR35IjA4ao01Boi+oYPQoPRb
REcuFZ5rZSmTmYwhQ4jEl0A9u2xLHBL4b0Al2s1RvH+RIyBm6oci2aerb4oGNDto
OUx9jJb5LtX8m00rSADiG8lNOXaftwZeg8UgIi60UAtoknwHJzMGUwGPFaepndOL
cWDWOQM3G0deqsbLiILXR2cHN0Ld07I5aRytUCZcdEubbwCms1BL/TuQfAMBhgUe
7rFIHwvlH3ejvw4NzWd71UnG/TeTuH0ow290K9TXZSleaXErpMZSHva86EK/DaK3
114V1djrKXHb2JaHOW9y2ArKnDycWWwjywgS7jpZgbzX89UYqtDao9v5a+MbLyKD
HbGIc8EvnH3QIh5D2BTYIQyo84uIXtKot0+tbJkhul+EbgVP9QOBzlpJ5hiL2AR0
B7CF2FmohNMp6IpDEjp+okTF+E6y4ca9VMi99o2jLEwC3A9Ra2O7D0a/4LskNTgl
ueN1w3bFigtf/8oc2umjhYqwCACNB1qPXRCQ23KKpj0WzpXd8bSbK8oTfZ2Hh0rw
k78HEoqPNrVpjJ5HxQd+Tt5e6ku83vXhiLMxIvxAWA0ItUx8ZDgwcQTI6i+hDBQu
N3yPXWU1LJaozV/YMkIeMPxJwBx36Vlx9CS+G6s2+NIUnVJndbLH0P2xwJ5gRM2d
1N4dLna09IFpei6aOha26dCOc53qysPPX9qKYCaNj64s2GV367cpURpIpTMFjDbC
Wo6yFHdnvyDLHQlthyaqtDQTUasQxF/bpRekQ6kR8YP814do53Rg7Ep0sdZjo4Dz
Mx9q8wUrOOTOf/OS+PfiItZ3BbiHXDFj3NP4DPXLwILIFSPVhYPKPOZuSma5iMnM
Tu1tLl7pEmL6HVnMFjRSqBolQqe3Vb6sxH/82LJXl5dL6UyyASYJoUfDtMwPMmsd
MGTVJzQPoThCvZnVknScMBi7arq8zJMfh18P54qXhGwg3vdXmahUlZuKhNxKlb3u
8Nv0l+T8rCGzgN9XSkJRG+R408aoUPZWP99X3FdsTtNeDjP5MBVxYZn1ml8x/zvD
YBbDE4r/ZKlWLr4MAiPODroKxykIqJGbGzyAIQy+a6m5KYwoXlao13juWIcvsALS
9hdOLHcAkL5AOXnzjVIbMBavW6bt33pSkQ+v6Z+VhnjAswjF+B1FBwWhb+/rqeB2
3lsqlR4a77n4K8Ep37aBQWBLpMFxyOXJhh7Wn/5Y3WSwe1KMyXvRouJrwT8xj79M
WywIKQnD1wisMlND8rnl94CQ1EAqxQ4j/Gs+DA/3f3TYTJNZpO9xzMFGgQi/Cm1Y
mRiLFwBimGz0PRBo+5V3XlppkvKLaUwrsZ0AN7romoup22OnZMQST2AvTWWq1e7R
G35ypnEvSXOodB4NTAZS7bg8qM8tgm8UEbGh4LAUhkuw8MFPamDk2CZ0Upo9UMNj
Ve/JQujYskS4+UUz4lWFw/wBfR4GWbYzPzb/TOSnxYibfkRjQlPzsc7Yyj/pyRJd
RgKcDHth5qRaTDf4aR88GWMy+18Yoa8++ic2vBg0wkJFcN+Oz2hRYBu0l83UtcEZ
OktSNqNKnSiSVjbqKxVSatVEh9jaLtawauqlQe+cxlngAkQya3KboAdPXB3NmZ+h
OosVElLsby170o275qZdUm40b7qJJHSVwQTZn1od46ImdNsk3TXYCJhRgLjl6feU
zFNUFKu4aHjidlH5YoELw8R0sQVizrZpwnIYZ8I4imDG/lES6vScOvFUQQdF5FRE
dzAQmFDevFmV64q/lvfI9lgxm4E7xeMgiLS18S50q13/jJe59/Ujgu0Xn6iEsYEx
oLlH12TTvewN7NNpPgap99AIEhAwthEfemPLIuJQ2BNPydjovaBcMVFne+le8fwV
cuPECAc12ctoXDB1+gZNchm0QKut5cC6SCEPjn0hXj4QtILtmruksXDpJqZggxc7
FdwvKaaR/UFw9bSWB+E8VVS5BdBt26pVJJ9gwVwqLXs46Hijp3oLFRjfvR400qM3
QgE7+L64wbTKFHzEuhy9mlMaEf9t2y9jr/FOaembupyegstJA4CFnqy948UBYp6z
vYei8ERMUPrQyvkY3Jay8FkNZ2Py042PB9Bg4tqu1W1H7bIioYVFH/QkZ85XygqJ
wu776oKuxdc5vFFEe3IN/MVFT20VrB/tHQYhcUE8GGOlPYU4cTWvmWPvHX465/nb
/N9fqC29M+ov7nTycPfktFQ8PJhkXlV+cef9wmlOhAFVvYexodRo1L7r/C8CnEFf
mbgIzi1rA8FelTdRbEGTe1RMvncCeqFqwzoj+ynIuVtVuNVUFkzg8WzW2Bulrr0t
LalFaiPhUcOmstWkuUca2ec7JHzmpDQSPGjvlII+UOCtSlr63wRyIQp6h+cbFpxM
qFRJUijD32JBxGefr6AwKA1+CBi4oz6lGjGO5Ft4YMrCoTUhElXq3WYvFxLMSbKV
cgCvDdLJV4sXCYvv182Qv0rDjUVlO+r1Pjf7gFzHQSFRczHnq6S3UwfEMoRazOxk
pz/TJ+cGJMTM0k6jTZqX1GiuBwOlcfsEW7isKsJ8Y0OhRCoD3EcFob5SLKjfoddb
ZYZbPRp8AnZhNRnvtgzYlkDR3tITBf0LwveCiVsG84sWi5mA80akZN/bKDrKfuDt
OrVvF9CA9iBP/ppsK8zsJWY35/d24g91+cfMJuWU7EZcHOjrL2FElvcOTsMRgD8e
bCXD/KC2mjApt0cA9ZQQM9qxoLr5TpP+LqZpvsCnKxypumjPeYQWvWumIDSxFHo9
3lr7m9A1PVnWrI62OkCVv9mv1e/0AMP3h7/jVk3TWwiZh5QTEcTt+one8PbZraCL
ToN9dt+cVfb6oaaak9NKSdiXq9GuUdBAHGAm3/oopPRNQB9tGtLGCAOaz5ssRBDX
OU5XUOcyqcxu8ajnN4OkSUkqW/kfjFk8/bdueHaDvZwTIDCMmgjx1MZUeOpAUg3M
SeJ4TK6XvaqzFI80aa4fLlUUNw1viudHttnodifvMaXDzzCMh9KgwxdEklfPY5rS
NjX7E6NhK6gltWuRflGPZI9kf6n/F9N+Me/+L0ImoBAp7414rqzhm/2bHzkZUQGF
qIY2P6UzI56OXkshnWhV6JiX53WWAxQvlCKGywPfL99s7hKKmQPth2dKW+pT1aKw
voBn5OV64Jjml5f5Ea59jKfMQHZSvHxsGlj25zfm0Pr8PocFJgSlAa/EeyN9H7Hz
94YkZy6T6BnNGCAgnB0gWu0C5/0mWz0gAN6AVPoiiL4czU6a4N4yncmLoL4PhNYW
I0yj8bfIEInU2vKQ9/c2xvrQ8vJfRVmF8NE0KZHb2TsU6Xvj4tV5Mf+dY4Iny73d
nCk5KCMJLtYDnoiL8yKQZwJXgmblqPfjashCPbbLvuRjLEENuU7tmsjXmE51I5BT
1IUuNPeb8e7M25A+ZdyB1j4jYzS1XVEv9NkwV+hiN6uAKcvEwQL0n6ldlbq1xR8S
/7Khg7/AOJWHmVOYo101T9I/OQMt2EzPVXJK/GBEz+AeoYHZ3FB3t9uLJMZV+zz9
0zIT0ns4FcLREbUy+ycpPtqsKbq1pe9wsUGQtviw+CXAv5Otiff+WTExxfe3u0ti
GQG1Tg7tS2iEw0mlwlsiGBQFDmBTV4ifPaRp9ZS5IaBgHfpg9GKkXSwAjjPcsRSO
IlLTpcA9xmoCOx2EXZwX/9nxmSxShPk/DSwhOr1IW18o71OJfbkJMqtYBeUefO+3
0+17mJtZnvjHMIjZZLQNyjN/6OTbkLkflCkzJ8Wmc+igjOeCFAp/4Su15x/1/bH0
4nDVbWHTCJgVIz3DORimUC7yTI8iONHtDQGgjNVEUi8S4s/GwlUExLXlkZUPkKV9
+f8W0sZdSI0tZoZzmldSEE1qGBnWID3p98VHBvVr0G8YQBdifP5esvkS8HLZYMYf
B0xKJJaxd8eykUUmUuiGaiwSJ7UGXsw1Kan7Ct0HQpBJlQYT3kg9eoepr5zwlg4a
V4fkYFsU5QSXwpUuL/ECVJHiqAxyA+5mM2JVBEL3jqV5oBy8BGeC7XB/Z8NhTAJT
kzxST8tNrx1Yg6mj2FLdov3fpKvailaRMVctpljg69D17rRstuqTh15mJpm4GJDU
geiyhVRNOpUxxVPDGJGccVw9/2tjx929Rmy9W1PN4JlLNlYqRsJ35FxuFr2LtYJV
CkOilClqPOtCOQOFooKZ00TF/j8lD66voD759MnhBEMtWbHlUbE8VXE4LonKy+lR
FPb20sxOaC0WXxh4yn7DOXiWxHpAsALpIhXTgPqsHJ6Z4u+kCaKYKDL7UBunVFH6
4PSb44sMNbxEMDTc0J7N2SGkPD56wTd2GKTJ92Fstq590CZDwiySzeiNS+yABQgw
4JbJ3viyamX+g+zI+U3X3B/3IBQmXARREglVZNHwLKNuOyVvpPEb+qpHeU4fVQZh
B4kK7DeVRzmv1swoUDbMZChJ8MAKxW19bvh96oxjI/Eh5bSjlY7azfjEdCEYX4N8
RRRcWUBpl0CYw2JZJnvbWQh1LW2Nh8gpO39j5AIvuSW5GShetTSYRdLPF7qpjmuR
deGznz7D6rF//s9qRwNMYZtOQzeTOnpoeCoe1oGMvrF+wP1uLN78TGceaz5RD0eh
P3aYVvaioGPgeARIqFFB2qnVGiWC5WN89ewvKgnEEPiJTycHXx43F1v+AhT/Rw73
Q5Jr4rGAxQHwce6ncOQum83N+qiTsVn+H7FC58go1233pxoJbBHrsyKgNu4Qq3bh
S/bIDdOWQ3JwcUNaRddVo869qCSSlSXw42qFOhOoPxUPRv74RAboavZAJnfuPhcJ
2fAxJCz5xJldOcz2bbMtKUaBn+CBSXPugWh6GhiijqMMNBJXpj1VKGBAKDa9cueP
HML2BY3mhHG/6Le3ol0An7csV8vC6YfOvmMbiraIxO9ni4JfMSCLEbt6sskqkXCm
dP1CKLVecmwnyUWguC5bnYSoc7DtHUYRXIH/ephlJUyDF7XU0rysj/kaXogVD80b
cqz2WtB1Sv/0wJwKeRDG9lSvHqDajBvP0WjBcmLO/6pKkoMr2oG7q2zUkegVkC9b
3Bd5hLerrvowBVB3u7ONV8vhjw7/ONUMB5hcCyUhOBmM/92A2ldyCuybw6nArvxf
wh+ZSfCtBa2hE9xnP1VH7kkxggZ3/yGPf9NTUW0Zh6PF5ZSSupK/d4gGm3XyWp47
gzslJ+Pg4o/7eCZyiVsudSLdc6R8EPJztJhXw78/ewqqp6oF2oipm2fm+/xi/4qR
PgRTkBPQ9DDeMYRfQh0Ij0Yh2//ewoHrUAJ7k6qLj7+JdHF49uXlTRmmH6E4cQHE
xYvgTOEfE4U8Pzp+I6a/zRapvDJI4Q6p2mv+EosU5dpMs43V4Tka5qi806jCGrxU
fmeESbGsXQcDw3FWrZ31m3FhFUiUltOiNBY4dBEFg6uTPlzWd9gn+QT/KoQdtrNn
7XTD9X4Q11AJkmcUkB0WsZDswCQHBXatTLndFYOrXQ9Hr0Zo5/sDQgE9aWGTx9V7
J59cnlKHzNbhq6Dg7Hmq3O4BrBs+3IE4A5adWm0jf5DmViY00FR/xZTer2ObPyES
tf3ddVnTtuo9wXZOkLSdY8UmroHcsvQ0JRaKU1pkceT73ac6FnGut3FT/SDnxplF
UaS7Wn+JbPHSvI7YaVDrcwd84a4Wj0ou0NZjAsIl9uTfT/0iGQaBx9i6K8ARxN4U
9185J0Wwxct2uxS2S1zQ77PZllTO3FGdt/6wFbKD3XLTKb3r+JwJzwnvqsQPfji0
wHSDhrpHKhNqwvmm3rsmgwePu0G3vbW0qPqCj6qNdUqGxpfJlfxj1wrUum5VeV8m
8sAyiR7/twBDML8Q5vdixCXXoolYrFuD2j7HBlk6tJghNrhPH1ybu5dG9luvDttJ
RciYhUa07T7irUxUIo19HgY1y2pw1EMj/AsRzjWQ22Bc5qtwC5d0Y+HxOLK+C4Mi
+NKMv/uNz96NVl7+SXiSLqupC4GST+44GHNVoZszEQVaQiA2yymwB/0ENFHdTqdm
UBROcfXk02kNjGBp3z8I8eacIi3S/4UUfAB2rpWPSKhhUiE3KsrlShQv4jKfP8pB
Mr/R8DaBJqJ9vC2iI03KyjVYG6C8MESsMIeou7IjTdVXxaomJ2gsHDVelv42VPFj
OL8hCjDRql7vXcY4sm8MqMa974kWDB3vejBWunBKEV31VUz7FaGQ1p+DXoHC7dRb
GJS+9z6jIDEb7/rFEkimHF4nqgfKCWulGb2NU9rnzyR00aTmlb8eFKg2wKDfDzT3
+4dxy5dzeymmai3jwtqAuu6Xl55kT78mqDRfwxlL9xI8iMQ2dktSGKxFG4RsdMKx
5E4wIVtqY8gRISdd7LeeFILlJIRFQg5kcpTjq5Z6cy9hxuZiFQhReZsE9tiRQv5u
2Ya/LJE2vFXFZlQ8VOU0cT5fdWT6Po44x36kei/k8eIGc+MpNvC6VTRd+OehkWSp
FXdD7HEGk4Ta4j53ilenaoRyrX0JHYgTOngCbJBiivBj56QTLcz0TWeENKInueCa
JSnbZJlw29O+ycidpGJVk08oswirwjua7NYLGyz4vU5v7w+EZ1qx3+yFGYmBb30d
w/1Ncz3yyttLQZJI3/1yRWrXph67DBAMCy4+Hl62QSf8rkzj4Vh7naHeyRvueM7J
fftIGTjKoev0vxCdiUCUV1qRCBiCXrtLysV86hqE8T4Ijrj94N2HkcxRrNeLYWOs
DsnX0Qo2e71HTQT3w6uvsdJ/GeFopT93rHck1qd1Fnn8BSP6AWFXPd14Fk7vL7Jq
vNLe15SSRpasE3EJ0T19wkoEsE8Bu3eBsxj403pjOm4hDydNMGRwILHn5HYIJitf
BmSGt4yTb6nKvq/sAzaS/y3Xn2oljXID/mliaUJ6N8aN1Hxl3FcHbo5HznsgX2np
wchxe2GTlKwrdTf05Rp0BqXMdW4Dds2A9TacQNtQeXBJJRFauwEUE25TCbXo7XQ0
h15aDmEzlSodoo7F+Jdl+OCprqv0JE1hzTTnBKLUYfolZN1RaRItCjLeEDRhYE1w
p9GKcShJCTlJ46eM3tNktj6pZpjDzRRKqy3SnB+/IkzzP+gFB6zq8Uo4ZBU0K0p9
14XLxz6zDeqWh0jJnngYUVXOdlupS47uwQDpTDIdJpkW9r9rTPD3HJhxBPs8UoL1
hnqFUDEq1qaOGPt3MrUbYhhP8S6UQLII5IbzeG5s2o2ZW1BPX/1YljV44BaWFLl+
PryY/ZfrHp6Hv1gF77uXrdxAAugMi2dDUQVOcBnZDxTptVkJmiOJsm6QA/uVDOr0
rNj4jxHH4hm7PcvZeSQ2G25TsR3CvVeyn1uJpepYqFn6E4iZ+iMS+FflpMMZHC4N
OhkI0EFvVeyJCna3rNAy7zOVwQouomkhyZrFYeKLuXK0m2UupAh+G4HJkiSDhPP6
WhgtvomFDc71odh7d/3vbO2I+Xaw79lLajBzsVw2ZBiW7cw06IM7bfBUGNqzpyN4
Mzyuw6LmawrGeItLxtzCBPIfIoB2ozLld/l5HdlFEtaaTsnYBdFP4pbyAcCg+8xU
BC/1I3aOG4CujNOkLkQVNyogVuqFKLLYjdZJR4Uc3CS3CmvjiYIrySVuGS6dcQ/4
tU6FbpSdOhnamQdPSt00kl99ymVpV/9iDj0fsmlGPXjDWsFIoJuWESTedxJ2smwm
Uok5HIzIURVwEInSQ1uCt1/benHLFQcPFUOD2v2IUEURNt5uR7/8bUAhZm6qnv9Z
oCJw3FX4MhClfHaC6gFXkhEJDrWXfXeXI/WDcYDR7ZiD5/wx3We1ENt1tuWN5zR3
juCaVn1y3fXXHzXwfUxmv/p9sXJXHQg16dDHDFYiQ4WTs09thRfpN/9CLYc+MtV8
aKdLu5DsVoDR7x4oV48j8n812+VkM8sG8uEiv4d/z6NDE8/lrqbnpsjLQYUTKA9p
6umUAwmNCkZZVajXLlwA9XXWxp90h/0+ai4o/C1DxH6/i84oIgxHHrG05xZIMMiI
5cLP+F1Z7NWgYmWJNyaMVrjMqdmDjyPt8ZRhGusCMeScKuj2vp9sqKNFk/0PZ5NE
FPDpH+ahs+iSvIZ7ChzSgUJaFh58xP7Ul4ZS8K9xbhZfflR9LQ2lsNmD2V73rabq
Q762C/gjIsqvVdMZE9pg3xkJiVwjIdNE0e6gwBm0i+bHj0LhHzOT4hSR1IsOMKQM
2rA3yt/kU7yIYxZCltDLIhawQuHdZZzY2OouooC1Fv8WPjVENSTplLWD9sDiexTN
5Guh9lqWiOwMQxheTWGTtZrJOK5PLVTaD73dx3b+6aDkWmElZ1dCbtpBqHueVzIN
WEiyNT98A4QLBF2Ca108hSUxPDeZeGbsT3slOeBGb4heCdp5AuThrt9sXNg9xQbP
P8owfcjE9Jec37H/bQ306yRszmQgG9aD/ti8j8oHkkheYEFfT1q54gDCIbd3FTS1
bzNWx9Ri7THa2PERIJUVFuzvIxJqlfe18wnr+QBaX7fbWQmpEU+JCuYfqg2jAUZ1
uvwyD3raeCXEk7XGvbVZPMnWYf8/YLAuDsxQLzexCSYma16GLZYgRTCWXkEtjWEJ
U9+eEC4vGluGPWVaLU0X9z5FIZKE3rhByaFtTKtUvgh6I0dsKADK6TPTfD9TgwnX
RRXMaotz76sqiiePUUSQXZuX5CZdHieO39rSGNVlV19iNiVWgCJVpL7v3Roa/4ug
WbtavMs+tJvjaJ0WxX4V+Bk4DawAqrqZfyogQOJT3XuXrwNPTEomxRJe4wSdRJyk
dWMiFIkO8SLBpWXtIJ+LVaL3OdqvFBZQCIE83f+VE33ILmNfIBrd0UGujaZVcUTu
nzrJSf4NrDBMMe20co9BUcvhXI7Bn+4eFv5vutAw+6hFzBpTNkkRdugTwQJ2jaoB
+voQDFkKYEZMyNeG6fisQpJUG18FRd3SvCuBGhbZKg5c51BKYyqV/lkNXsy+J4iA
MwgC07Nn66jjqenO9XkZocb0peT/1HIgyGcfCjGQivoB1+vRqpQAI03rY/7dU5Be
+SKBNx9AkFwgB+UwCha6bO+7h0C8EkaD94KvwqifWZgymEM5ct324gV3aI2+n0uU
aEc/fDFi42OPuqK6YAxoJ7vz1vIqZH373LUGQVriprKD38mi8oV14rVRX4CdQLOy
3DKwt7hTqNi6nUCndNvT5PatxL5ueS5THKxKD2Uvhu1JgTaSuGXxwOxFThb7TwYR
RxvlNXF81ZyzObXs7fhx39DOONZQk1jGFvop9cYfixJLJIMHGREyIEhXVFmK4qvS
3fcUmjBG3PxybPVLiOm1SmTLCPa0bo6nz1KsBKbGGalAXG7Y1yNkX2j9JiWahujt
RktaYIE42upnHaEhQiMgF3qXcKK196b0Xf/p5IxLPEwsIlYH+i/l8pbwjEmYegpe
BFfkuQPn+xlq4lbly/acr4W5WohLumo4GQ7uiVbruVL9KzGfE0jZy23AIbzl+JRs
OBflMog/Zs7otGPgXO21SPnsepU9C6uD/D7mRSnbFtcg6NzKPNcBNt4MXwb8B4r3
Rz3ZVDxKiLphxuLvwcKL9Yk2Bb/RnEbgtxPD/BqD1zT7sVtM39E+pBNmQimEizNe
vudTE+6cp7ScvVbxQw54Mr8uV1Mh8AFrtytLBEKg5cDtKlFnI1ryz3GMBoOIwaWW
KT1ATKMakU4O3t/nxA33c33ycWj9cFIiW3hsZkvrRfqEdx9Vcj7MZ0/QY/Qi81yW
m7BYk+/Sey4czdes1IgxINToQRULb6IHgpFqpmqyn66j2ThVMmLoK1HAECCNzQzs
7QHSTtVlUr3H4XT1qNNOFjRhVzmICzV+CLpPyHfZxUFxYytWn0l6Tkh6f4QS+xbL
gsKO3+ppRBUQ6yLJ+9XJWAYLJ2BlQZQIy/6UyZSaEE7aw81XhXPEhvIWkDKldB2B
OOttOn65DMX2QHtbVQWzwarlP5Wpq8yC4BQ0Z6qIfdA8kY+M92qYQa16xgNZhkD4
U79SrmFHY0roBPmLS8ku8bCsevf5+EH/vj7X54hxiQwHKE49HaB4FZoua9eEwClL
IAN9HhVtauT3Br963IwUulq+f/BPqOLtUGWHmdJDjxRae3gf4oYMbw0pwRmImbLU
e4J1vwq0f0kv9HUlG+hchnXzCnPVg2nk6Neihl0YX2BoMUTKmCeoU756+MEn+K0Y
4D05cgINdyzmiZk4CA2MBrEfPERiUzqfu2WFysi84xpcgqUPohSGCS/PF7Mehg6r
A4meDoi6QMF/Ijtn5mHogvQbEIhtirSRrVA5TF4tptUq4tHeulODzmUzeY0ZcO/z
kxd9sj1Qpf6bKHc++xxT9/1+Fm/W25LxPNSd0FUMw7sAcUgueUVyhQFJB5R2Qrs/
bsFn8zA/QYGpft1z6tpPB5QSwBdJO9KrMaaaG+clR8+Q0MHmp2afsSIOEbY96lCE
4LmGyzj8SW+TtdXKRaE89L1a/7IJTR728iCrElN4q4MDGplV+vwZVQmybJ/aAUFc
yJCxpWkDJSMkbBApqct5OPuHxN4OqgnryFWuE0s+2/XDTx8/nzONd+xIXmE7F2Op
Yp4GwPi4cMxZiN8n/82UUCwr98ppqlBvmxrbbLXbv+9F9Z0X9eSVk88Fl0qFn3wI
wYtLaXKW/Js6/ALmeQSjJV8/grgfHmMFQvvf1YAFWAZ6gpIWAHvMHdSo51P5Xsfh
dBfPKUyHtS+JQiyXh6047RnMirfx4y1gQ7BZv+aNRVVH+jpAqYCUC+bSkofHqUIJ
ZzXoMSfdcBWkH+UhDSlAI9t0AwW2u1Au2IyomO/xCfWOdKwYKDFABfN421w+H4eR
qSDaG/IdRkXi8GTYDZiukWduQbsAYtVbPE0jLlQj4aEO+yHfD1XUokECzdoNtKHV
01OZe20P2FZNWJhIXJAlXfGaCDXckltxGWOv2XrQm9bSQlhep80E11scRcY0+jQs
g1FpVtUOju9H/mjEd1Y5iOp/QtAIUrcerWZjyZ16QU61iq5ApMJObsLEjSDFnklw
TQ0oJJ4SdF+sys9RQrtgFmlv7p//an1BpB9ObDBVnJJvsssLUnUlhWDMQKCybb/k
nOOrvHRdg8blHf1fyAbHqo92a24QGQtRlIEHjmC7HXfkX5OnyxlOREoODwLvsr5Z
4SzLVjcGj0rEJS39aw+4NrIWi13yUQqUfGH0cVJYVQZRlZ6wsGmHEPJxfmPTGJPr
XhlwLGrNApqFHpH36O3ILvM+LNOJRzTciEPKwvzp7cBgvVILTfeCnFNfMHkXJuHd
41UXYY68u9N2r8zWK0LNhldeUG9HlasgTrRuVUcXNkru87Adt0w3805x8w2wPDQD
wKEF26dpfzpsbi1rp1pShf8KBB+rGuHER/OqQVUl7KXhEZ1N5pRxiCtVDfGzrNuM
b+7GousLvnpTrXf0Ltlsyyg+2JlCjKptpQRUPGwd2AcP0oQgxLzWzMFz6GdoEYyu
dbyj0lSXiUVqBdlukS0n+tmntuSroJhLmjQ8MlaLVEX0TjAHycRxZmBCa9UvV1cA
IAL2t+B79BEEPYlFDK536RqL2DnZjku3BNs3yQH7Nt60jaFAS8EsWCrNTpS0Rr9E
WYBl1CvgxkgPFd/h6HP/6TJbY24/SeK4qrT94RjDx7MZDwPeZAkSsc8INfJICLhy
n5mIcsYgK/gVP0HL4dRp6T5L4/6PTJcrQg5b6Oj1o+rAsvhFUNSKrcbu/iD8OYNV
jFZgBRCAsKwCGJxrEH/HiDp3XvcJQcOWBLNchcvUPS4vRPyea4Ymd1avLCaYHliz
kaGHzqt7HyWR9NTFjNdQDAV1EACF5OVDYKLk/FGhzaQ0lFnXWWjRR/N0ZUoN++JZ
VZ/wKAr+tAD+3gkGeluicRF5DLN+yF4wsgRsEDSP9EYXcMHSCtKSFHkWs8RmhQFP
tiVnGSrZm6R4rGsQJLtS5G8Zph6pbWFT0sEVbJ7iEx/Tt9DK3CjP63c3tSeKqti/
sGGwwHPrElZET6INp+00OnDaSlJhjWVpgNbOhH1o/B+LkLk1v+cf8W1XSezX99cD
uAXOTXes/UXtNdiY/F4jz2cH7P74bj5oogdvp3fCNoR7wVA1/7Ur2wEhr+YRbsXs
xOnNNcPkgJegBi1a63k4HWLxeJW2jUSx+WU0i9zCnfWSs7DG8JNs6FUayAiK3u8M
hyNvk1HvSZTKCGH2FEldlpkN+3k0ubuLsIZtLbiEbRPTkUa2pV/E3gJoKJd3jwUj
h/qRN4Gyfs/cwy1QV5OgoQTmduIs/xyM6FNZizcEquTruh7RBd5TLHq+GSsBuFhU
qcvr+AJsxz3+F//gYh2+4aqTzf83RDy+C2bQpo2zzRm1W/Gk9APEVQoh2+cbmg2B
RCA144W/PXFkOTtS8TrpkeQwwy+vK9973ZE15HKTESwd0ywAMKEcLo6x9vM9G/FC
or/p0bY3r5Cd/UnsjcWfKAuXh03hhai+Qf7ukS7pdkFfwmAM1MtbXW4PthprcG3F
O6xTe0L31eUmUiH7wIcO57Ak6F+cln8Ef64CXj/jOiEFc29k/ewF525olKwJ/4aR
WkoyGWRLQcPOu7wQQdmzhkP4a9m748RLO0tPP8kziMyDDY2Yl0Y6E/B8AMW5pUgi
CgiEPH53zd2/4iZ8JeXNdDnyUaZb3wdUP3F2UOPLdb3HLK1mlGM/Fa3PHB7EyF8t
Nzi0iiEqVI/Cu3qjkFlwbtIY7SiZdSIGKPHhe+gKM2U18gL+ZK7w8Ub/2cZhlKnw
09PBtEixmb64Ygy3LXxkUFCgOroLB+LaLyL0433fJuMnBPLkfKtCHhhngYPjW2VL
cjedKNmY1jSAr0L+KVdBVQRZEpkH3lYgv02DlmHsIqVg+UN7vDVcxcffAZx9nI9R
5Ib3q3jy9V8hRVu++OTlC48Ku9P4cuQMqFJaZdurW2g+ADPTC9yPTmk+m+3iImhD
LNDhr+nmAlrwmy1GqgJJEUdUR1dYf5meGifpzZqlgqYE6mrrE6QQ0tFz1j2pr2/7
tEwR6KJMmoY5PgH3xMyntmrytZh5DVSLt6QGoefd3IUabZog+7ELuWtKShW2tSym
PX6FYboNcsfiDzh/6CjV4F5OEJ/ZKxepYwEnicXfmJbIO06cz83HkyAdkl1NhkI6
YZ2jmedcD7NeEC7sOkje96+8+eQkN+roqpPRmhRe/IoeOzcC41Xtpss4uiQdXP2d
Oea88GJJj4dd8XMh+0DlI2SWaHXsxN+tPaXYVfZuQhOOyY/T2I1uhi+RfWZsNMsV
FSQ2SxrdDvDmZV1p7hHiRbB9vyEK9O4M5o4ynM5nJ427aaQkB8KkvkaFz4HxEunD
JZclwou6bORv78tz9Na3wX0aKAp3JoYGpvA09cSumvxhUd4yuJnpIL4FDWGVTP9a
7C/habXrW2tq+rTq22IFaf8aVyEs2i1EHGEgjBqFysDRPbmNO8O0dfF1N+xt6sCh
WFgCpjz6XQ8WkSAQqG2DRMcryTqfCQQJAIZoG9YiHeY6bJB+q48oXT7MOuH+WQok
hLWVR8HoesULgpTz0bUQa1g016sph6lmI9/baukomLNBDyG94FdZsCCprOS1CZvQ
95BNfbD5m0NH21pgLMBhu0849CD9t1ruStHbR2Q/hetNO3V6nfaZxQuiAgeekhPP
m7mo+QMXps/WwK6NbBvKmBAkkFHSBb5pr79RGRcs5o2v1iMq0nbFcXM9mMYKqkBp
gDv/9KEJcENnGc/TiWjbs7XLAiyD6o9tGt2G9Tkm7FMyPttoyNilj1lmtVFGlgFL
Z2a7DRmenggLMsclXsfa1ntSEpcOYH45Z35s1ibyRFcaBpMnmApg4Du+OyqMI0Od
JJQ58HQd/TQDw0GyiC4AY6NWrb204rJDlLn/Jxi+d3mBZEwcUDSSCPQ8USm+7aUm
4i8cyXtS1zq6IxIbLYW3ajbKo81H1Uaug5nQDtagLqq9s/lGS513ImoBLKacbZGp
6vhdElpDP0SpjE/gWAal/dUaPLt+d76lo5kCYOtnhsl52xnjcfhQaADYwQt7fdUN
BWEg6h8kHrO5wO7eUWHrD16brN2x8UognNvSbvLJw+/kEvIETJ5hNCuQaVe0vyLo
lJrCvlP0cifYUq89ttqXBh2qJpXcIhA79fTYbo6Vz2x4WJjPgrUQiyorWGla3GYb
Buo8KUZfpj4CA+Eth7aMBUO+W0N3bOVNDzKq/omEPW9qMpxMVJY+//sid1XUxoG6
b/+nAxxF7acMgCjuc39WmJoaOgKMpQzJGz3R8yiEYEof7IAI1MrjLqUUdee6V1Cu
YIAJNlLHrkzyt4H0a3oqepTZf96OnyEOGJDLkfxjcl+RpdRscXKRsSDEQiYoDk6w
+QuT5jGQAuPw2VZj0YTbiQyIvMnIaJatm3wf4UEBIBuyIo7atk7GXfpAwk+QdGAj
nlqUWfN6AwkfxP6+Hhwg+GtXZDZgEU6jesmthsQfWq11jBN7WXB/H7Ak+q0XWLmu
rfUj3gGiTMQzrlPe0FgIh6RJ5XeerHcP208gkuOd/mJ7E1xS8CPgj0v4shzEHCsD
3f43vd1eONyNqebDUkGTeEbIidt3B2ZgxqVWhULtchWilIX+qZyOWkDOhzAzCDvz
HF/txO0dEUM9Yt2iux1X3BM4R44XUNNkYeX+U9yyLIVHjqkJUND+FaoLwx/w2OU9
G4FrZfb9sVK9kOF4PJKxS+2ZTaZb8HoAWriYWCmukwAmjMYr2W7hGEOSufrvMh74
ibN6IOsYXZxDp08EL6zYNW7SsLgILA/VYaXEi7lAC9OD+2XlDRDubl9BA3b5NfEf
wgYjn3dLJtuR9SxP53ahj7ZRNPm08lnGAgCeRQNbeOys5O8qHOrnHLpI9jm7FKDL
ObreIQBSXUIrJYgmNAsfzoC4hTVWNo/TJwJpmc+TM1F1QWdieitXJzbBzFjHYRP+
69207nX4Lti5ISgp4KadT6uv2ImK9HAs7NL2YwAz6o2Z6oa2x2+05WOgwtsenSCM
Ap1beomQgPnPdsXCI0HmI6XteChvlvFp60KdTyiHl9EaOZWD8cuT7CyPGFI4a2+3
2rFx7HF9+tzDozDtzBiSLlLeO15xrwsZsGQydWUItHeeMpdz68pM8fWbQPFAY5ha
oD74tdO433GfWU2zFV3svsP+fYBMDAEOwvkC3QSHScO/4z6BSFx7SBkGUjQ0cWf5
ZoW+on89+PzaHcnWTPOpuqZlgGsqJYKU+/8tHrKG77IoEFKW3hx3B6SrxcAKklMl
TaDwkT8EcJaFvLQ2y+G1NlSnajpEgREmONzFq85cl03+D2FVI7ls4VYjkgBe8kgN
4uLOktpSyvM3VC5rzf6VO+24IWH+eee0zCNNhCsSlt05mFunfhCOBUpRPfWXUNin
Wa1LbeYLqBOBS5usexSB6jOTP/rpYXAmkXEHJTkrUdnYln5vC2uikO4+OhYINeeo
eKxOKoZ1OIgufqlIEvSDoDUEZPu5YUreqmnQSee5fBdP68Cx6VcB3FjBJrNl0KMj
U1pTFaBtAAdMTsYZfZRWux2wKu0Ber78n+uE4YzKUTvSeD0ki7TBv9JvSyBuaSSA
KHjYs8M/KFxQU5m89Xqh8W1awAkkFdGHDv7boT2CB6HmEW75k+vdWpgYwlcRKIok
1HZLks8PY/JqzTPB2xGzgtWOIf9bemGy4n/6XD5j3IGMFa0+L26mQjwczIz4/jRv
s4lflcStoNcRKOh31j2HYCbFhyaRUQDNidGlzoT2OyrsjYgKJ8Hx5Jan82VpBUlR
g/ht1hnDqfb1mS6q3QassV29Sk1v2dY4NCpCTi3cHMFpfKylpaxuex37js0M10q1
T5J9HJ0wFAeSMMqq9EhZAlPCXlzrO3LLz5OIRIjyldixxA6994/1FShBfprT67dr
ttzJNRLSODvnAz55Z7uu7pAfXPNw8DU2Rc6H61kzOxmbe/ohLyCVnneQYy+9Z1oS
TBD6WwFdFEpEtGUaDhUURknTtHIJzsmyg5+D7WamXbq1DLSVFuU0Boyh3BjdsYKt
S3jdwHfgYRR9WVL3lGWMVFs+qeA3H6a+K/DBF3wf7gZaNj2h1KVnrkA8smTRjMeO
3QKnxRfq6W0pcZOCkS0srGEnIlxxsaRu282dvmTtvnVL6h2Zi8eB6zz0DMlxHFrQ
I0iAVFta2E5TB4ecXnUHpfixjsnRY7TErF3ynq9vwLlHeBJsxAOioxV2cpeUN0gf
eyXrBVKKfQ+GzPNoHycItYK2/T7QjmHupkzoxE+By15RBte6MOYEU++n5/BUXQVh
/LsBlmsaOWJA/8ZqYHVAHtp5n88QtgF4W02Hn8Jogt+fQ9wohiBKpvaw7KtekEUc
1Tp1IWe1gyMHYBn2o7nTOl6/yObcyvqLH7WdNn6BpFHi4OH8Br5gHBTSDLTx5W3F
H3pB9ffdZ4Ux3o66PUR3q1JE3t40tyfxyxZRnepnnJtJtIDpsHWJA4B/8gUA04b8
c90mg6sMXwhwEGCH1mI/iREekkcef6KLcpdzW5Mdf+10p3Q1GQvNwDku1R3NspO4
dXFOiOhel9/ynC6dOeoNAND/BpSRUwh5LhgiaOaBsOqnqfsPonmV8abl2gFFcxXf
rJnLbuF5zSghQNvx5zC3HVhwGja+pk79xUZ2GACJlfivNvISIUABSkCnbWaj/RmT
+GA9CAH/CaWCFW+57Y5+dmA7QoLB0XbElLJwENHiPG1Tmf/YkY5XozqMKQYTGqJz
H78Hr9cOciJ9ni6w8C2PbhTvcM5/cv//v75OMhr7O0yoENJmuWEgk9hXd1UwksBG
ljTSZpuR4jMYlmXoPBaNM3Mki68dIxcyVeMNgOTrrHBnPxZrkUpJrE1rhwei//Yp
tw23TF6Fqy02rRWmKD9HujMqnsqSrYYn/vUxinExN7E2tmzpsyfkEG3iIrHZJ+G3
x6YLXyIkDO05pYUKCGxKXvAiwyeU1RFi8XbTk4rI8V/lfxTCZs0PnWnMDMV4BndD
lumhiGlC00vimkVScX2JDPU0Q/Jm+Ye4RUu7doiFD1Cul0cmTEYJcUjbj+Vwtv+Y
tR6GyvB0mhe2FBbiKggDbsVZdMbcw/oA6+jXrbaR+8fuR7caju0gasX5A5nrmKeH
Qy9MxbGAAXZZWMKYdKt3x0Tc7JPPay2hG4HvQZhW1uFPxwbjz20l2HKK9UfFEriy
I4k1wUCTdGrUlV+gKa6v8uOZGFLqHVEbJY46p5Pg1UrGid/TKAZFlPFxR8LlXv4O
KvpB9TR9cWbIvk0SGM1Qe/XpFwuMI8OJAWmnaQuXNzhh24jjnKYoi5mzutycITg7
UXcz4x+a1Yen7pOx2QCbasUlXHPspFOeopjkxeo4pSdKGqg0y1OkqgmO8dwpLE2P
haevTPUWq0q4f7EdnRKcgrJzK1lCIFXTcsg0urqaXzWFU6NtSU2wpRFDg9wSTetm
HPgGvxCbcPFEymayooGPG4H7V78eC1oT5vN5lLexBRE0c2pOKiLF4Y6lJnmSmXaJ
atEnBd0Ma8zUmp9ec3uL+68hkFYEFU73NqlOTeGriZV70D0HiXX15ZXT96FK6o3P
7xCbAS3lxB6G13PK3tr8Qglsg4Po/9WRGikGuZlp5m8v79GCf+YazhVh68boLabi
aAfpRreNV60gStaCwjKr+RfyJ/UNrpbxOelumytS5f8Y66Eydl84GRaWCUPxYUQz
Wo+hSLHKe8Ai630bJikugTLtZRQn/sSQ38OXT973RAGhHzdzqZb8q4oEINzwj4SM
ZKqHiwk9C6dbC1B5XfkUotKR4c/HpII/wYaYlh33ww7BAauiFvHe58sc1XAT2DTR
F0NphJP3dWIJrRyK3OMoWPeSlURolI6eeprz4CUOHX8FZJaAuNEV0URo43vL30jK
421FiqX+Cg6fxDzm9CfDF1BvcAAwmmPy29yYJHxAy+TSMRp3Ml/CX8xDwPuaGCJo
o65vPvlrcOO1am9RLyA3dPZiErvnWRk+W1mXG77Vmc4HXw9iSiP3K2136AL+339p
cWJ/n3gAnkjYvXuzz3nm0QPRhEgLtlWBjG+czXsOErv+ywKQeKyW0zjKxJ8c+Akp
kUQKaCV0zTa/qCElTElT4IW+cUbvBSTR9x2BOsDW8N2T5J8uSsJiNVzRn7rqRs+i
1mkO9j9iiMP96vvYD4JobJEYFWPXYibxVTmUJJ8XkIUhAJwdDpBWjUCQOEYI3t8K
dsArzLCnppcJYP7vCojQNVhQILvKS6sf1uoRAsHsqweKqNnbDRMrLD3RHLnaPfFj
ayWFkMNn+KKgoehSt7aEw1cNXKCJ93Qpr6g3FpH8+/NtTRcVlQbX1ZRR1mGHE7Up
8BY5WiRX6+sxk3OChcVw4B4xCKiCyi/MfZXNXOKKfgJNcrMIZo2+kyyY7D3+FP4v
Bf9+JlqiMbHtUsSlbAH2IPGkpjrgD4+QP/pE7piwEljN80dJQtKgIBMNWKH4F3fm
DKTphrU/WwVARJtbgDXMqGy1ESLNcPkVg17kiDS001tNNisLFqtlKldbLsjaEgXc
Aii4j2EChu0q/845FoRmJUx/aFR2oa4iSF03ZgBhT2g6l8s4yN3ybnA6k/YWpjxc
wRTDu/+ophT4+X7p5ijVMC9ks0T/85QUbCzCqnHInvaOIlEnimOltnRVPNDLHPDB
vAYIbLODGzw4IZxQSCT98WYc+/QE8hRYZD5J5ynEuUOfnVavYPqR/T2vHAESDeUN
k1Oytq5x08HxtL6wJ35zv1sONDeBu+wo+IIYv3cjZbXe2NnqKLTeDFZEXH5+2lbW
vjQ75hkOOSmC4nXYkw2YbOUyhZsdLXbumtVmyDDYNJuF8vwBW3S+LjYB6fjlQooE
QZwPowKN0no7Iu+T4uY4wJ/LSTUwH3LxkA1ALCXbjk6e2OeWc2gGHveGKjgauovi
qenDB8aMvCXrU8oEfbMP0uidoma6qmihy6ZHwQlMG2gsGy3A5JzbcuiBzGK24sWs
kGMcEyFnNGcoWlwlfVa1RQ3KjkZjuWHWWV6AVjMkYyRkYTtpnwe9UiK5qZhH0/kB
i6in0lihaMMM8RvkZLak0KqoZX2uS+xVSbOD95e3taoVD8/GhCwDirDSuIBiCi6+
CEXZZLdk9IFqsC4cqoWS84c7peODxag26mVoHk3bSFnW/y7rxZTqNIQcfZ/6JOFj
CY4HXB4Xl9q4FrgR8LH0V+FcNEckP6J9XXjNH+QIPDpw5D1XEPWuG0m9gunHDUDt
vYzWY0UhxbT3JEXoDyNxwVrNGT2aHidvDx+/GiPnBKdZQ8DQKRQANblmtZFi5KIG
Kh+rjgFixSn+/HlPyhlC44uFfRbc95a/TEJPO1jn6Uwk3AszmvQMqp25HuFXQv03
3osrrb+kOJJbkZ0WjPAT10hK2W1U8eFd85z5vG59QBu1lpfriNI80JzImlZf+G1Q
CoKWen4Fbwt9DcbSQ1G8Fsumb+M5EfdJMaHGlbfn6wQl+bZDT15K/B36IkfC21VI
7dsprF6OUC4xTTHUaqv7ZWGKwCwhCWb2xgh4KQayp7KyaALJoYo7MvSW/WDbUk7q
qY4NECUssGHMXJIY8wI4Wq0uX3z10DTSjIL/aXqlbwHuvNzue27CWqx2LAR6i2TJ
vnoMUCYFYYouyR/CqJn1EC9mkTV7jmsFI6TuQk2QydYGmRZZ2jUdfk3AObgnlj7M
C14fd5mjTgKHIcYQFcs0pgg9XWffQ2DtJAwTx6HZB00XrjqcWdJNOB4h8BLP1b2B
vOLlPfS/Oh4BYz0SMfKc4lXOzDQuM37sHYAwd3jlFBZnCr+HqecEjQgh1E+ZYQmg
Usyd86mJO5xghjjRq3T9eAdO90/hXttmRhew/5q/ateNMo0f1q5rd2N9nhO6JBi3
E+/rzTn4exBCdFd0hA3K1FBC9G4bI6uEjPFHx2xPZtv/JMA+ybfMcFVXJ8cK0y5d
v4SfU4vbvfRZ943QRVjakJusJ9bHt/aScQ9Jlns8rGAeIhaDlppsXhlzCv7L4Bg1
FSx0FDfHm7N3TH27H9QLKVnYUIRrmaoG6Ew452ad6R5Y2rtJHfBAHUKPtn9tefvk
0ZwhoxZVv6QuvW6gVfYMGMGPLJC1vRTVHcjuZ4Iwcqdt6aM/XTbw2EECQCOwMKLQ
1z7wzPKWJedw9tFV17cUSY1Ve8hOve2R8ou0mBCK0G3XJQ1ToH3O7+M7oGBIDjYr
bDD4nY3LNFHTlYUpTR6bMUHQVmSI4LusIQ0+WkENrHvVPI50FyKcQ0KKSXxDDsqX
8rTE4L/TpJZfOutfBPwVNgub6PmgqaC8B0FkffxHCQhpWE7WypOmHKK4Mdk9c8Rd
yY23M+QgyreTGWUNrqiPGy/GeCSKK7OkLP9o/LSYVXCJY1MCsCBG0xVtGzhdaWzG
i2D/TJPtqZNWXB9jXY4v7kbXCe20g92N2Hj9aZz8+ZwcM3NI04KQNYxQYPjnLz6L
OY+TdLieA/rY2PR7dAZtXLXmHyzFBfWDW8XaN/Fo58yg7IRXwkN7j83bCxsGn6xr
JvqdjwhJ0gFnuMCMQYp/tdZzt94jbgWmJ3u+Ji7fpd2ZDal1cEAveXBi2wMyga6s
yGL8+W9C0EyZvZ9jL9OCVHYc4MZDrnHj2vhGa0lpFedxc52T9fjgRqPNtJWjxlN1
el0XnbEYzTeVX94ANQG7I4XwhZUP77Nlf6qO+yIL/WJRYwB12LW9UIIKlG92gp7U
Oqrr3h5H21SuzMcypeBqW9lQ5UUYJ2o9C+mwWfd+GsXXJey4WfNHErELjaPPx+Fw
6Lpx91DPKIyHHh5h3OOJ7ENJ3ieDR6bdITPWdEoXhjsNHFX486FF4I01HgvqjjnB
EZXxioGcORul19JMtc/l5nDyGzPW2lBW+QnfnjrsOZxTXmhhbm1E6vnoOfxYaCth
yGAV7O0LMBFoxfeO4IrrAvKBwjEFksKMZktTWIHntLKFUahwU8/NO+6B5SvProYr
WqQArluejIudBOAPJQgDQg40TEDdoK81/VxjUqoOHW5SjAA9X6QtbiSLk8D8i1ot
59cRXqiyje9Pyfi8On36D5vIgfGPjNsEkB7DWOyyRTCVZVXj8T6Z06cIgb3DwVxy
/4HKdKo7Mw9mkGjQ97H3i5TNAqGM/57mZjkxb9lAACqkzKc4RCNXMzYNMh7UReVZ
5E+2iHM43a4Tqfsxh9Om1arNV8vDncIVXzhs96AOJnNxSWW8IYFLqlZSKlAM5k/J
HiA30f3aS0BetDvtELqeruUcsYu7hRTEl6X7CQWdBvsWPefnKj+5GwGnyFOnX9Ql
yyg1hODvRcHDlqYR+AVJOoGQrEVFMPqLcDvnAoVDtaqTjnHChstLFQdfMlZak0tz
PTqjWHQx1SVktjBbDrpzxErabF89XkqR9ifaX9XrzzkAzyl+TTriCQKo/wn525p6
q0iMUnFL7SoOSqJIeDhij94H/X2Fyj+5xjbvgGulxtC+UzDyFASHDDZWNIBtAJmy
CsH2IfHZittIrU4fj5mEoDvOBH612zvJ7KVw9JXSuQ5R/D//jAP9C22K7ZnzcS0E
ERmZkyg4P//3jqDtWxkwYFLqUZIaeENIb3iMgHRDTxnFehGI9iNxcX2SRyBvjSPC
y22HlIB767bBFFb6YRgvYocFkOfzBBe7IqwepUdP5+IStTqTXsfAcLYtRf5EUMUa
X1Kml8KiGC1pt2sozTpAQXYs0L/F2eqYZSEHhWzSQ3iA+LRnHGFbjFCR08uiEFfi
s18JOqmhe0txo33LHAN5YJZaa+uJVST1+yR64fAohbicNpT5ip2yOeOEvXxHrdxh
vzNfh4ZHDTmqgU6zEIZ3BVGDIan8kiHRc+Tje1G+HcfFNsH9Mo9LEOzohAdx0aqh
PIL0/7zSjyGju+49wdrtUlLgEf0ldEpB7CVvMkbWLLFsMlHhwwlmF3YbqXi2E7TO
h1+hEAnNNiXilVBOOiTAk98SPxjqr04+7E4d3tY2nr/lWU+/aAIQMfQpyGuMe9fL
3k20wLvVq2FMqgzvhSsyYwQoeIyUiLkZQ5fug4z78BY0VGoEtijXuhdMvoJYZ4pG
Q59l1GBf4t8jqU21Do7ktg==
`pragma protect end_protected
