// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
IRfwJBZCftMPPjpjqBuHyab/Y8k8+CM4IV52hfC1sWvJmyzdYU2XWk2jLFvr8wWhggQ5j99yRmUq
GLcRY502TFdc7G571dgcQ+z5EWl7mVxKssuEB2IFWV8cAR9VEfx3rR/eMDn6AWgbcbVuGzz8WMxR
tOdd/QAjTrQsoCS10ReR3QSKqUsUTzm1Qt6hYPep0kJivpaU/Nt5dHsRM0slvQMlQzDHWXdJRPX0
uQ6iBYuRfi9KK22Uz2ZE3IuRE13IjjmJ4N/NjYXv7aQ5MWwSVlJfC2VNclS55znGxCTtkUB4fnqb
UzJQc5gySsB5OGGBia9Y1gnw5CMTEbDI+nQgEg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
1380Sjlaz5Z2z9cf1WyjiPdZ574bfBEA4GaVuMWqMyllqMFzGrEiKWjXuDVpgNYHz1ajnXrQ4/v4
2VaSvLzyTjTIiKt7/mZG87xIxJEo5+K6WCAi8awihIORPIfWyJV4VGLxYTDWDNDRQXlUWUr/AotX
U0NXNBuaDG+y/HwSOks+lJuFYFV3U+y6Cf3HBwSHMA+sLDT/ZPndu8AzaGGokLiBdQFSS9jTBsHo
Kz6xwUQiX5SKryGCX4phkWklMCA6W9Dz6LIJo5WCxy2UJ0y+JAGKS9ysn92Ke9GFo2wQrppCnGVl
lWnG/87aSI0uEvsRyJV2W/NeCbgc2+pFZTZivpaJnxrSe//S4V5qIDFJNQLrjnp0pc43D35I7PPH
wMJ5jIDsj1Bad8pzGSTfghmGbJUucX5tfE8vOu8wWzOgj7fK9so3XO9NrGLQJXeR7hOEVDXD+hUJ
560pDZvcT1AlOw1/75AWJDMNud1ELPUjjKr5xoXmmPXBFqJZbTffIUpw1PWoAJbTS7oY5x9lbPuw
ksFtQZk4ojgboZd/Q89cLrSHz0K/YLOmkDXRyfXPympTFmVrHenTWJVvDa5EME/VxviINouwAT0m
KpjGrvgFzZjPkRrCEmi+DDThcpXQE4g4I/z/7jYLK/PJgEgSzEEvAgnYD1K2gOmzZ+8x7Meedv1T
7oW7BnPLrBcU1k7ndJWRUO0KbtnipKkfaGkezXome1dgLbvK5pWh0WiQ5N4suEpSWOpFuR5v0TzE
3px/hsvz1SGVzVnPCRM3RLbiJAai6t45K0XzxwOd7Ujd57ZIA0prery6Ez+3gWbZY/4YPQW2Y6t/
1skan82+j0nDhef2QYwAomxmaLOvi2MVu5M95/WqIVnEFAoKVmrRB+yJQ9vIvPYPAqd94jv7g3LJ
Q7kO4iGaUSsAaPhRSuu5ZrwTUjrnZdM++SSIO7H3y9VxCJMpp+BaRJKkxG9EqZF8+ywzaBasOhHX
ilhbQz40Ii7j8ULu3jaQJ0ujlQuiPciZcH31PCQAiZLah/QfZYPebqMnwtqluemCEUGnhug7VDx1
58OvfR/mfpJRD6L6JzHQSvQ/cl6tyJnfTQYEXxrKpi5zB3XQdvmWa9sq4XsqkILwsdGcqeTMK2Ky
lGZa3inG5SG81ndLuXGIRy+CipwUEbhrArHqkNiNMnbLaxvIGRTHcZ0aKdEFnWrnME2U4ATbVQtX
XmDcjhUSIlMktCq41VrXUEjUXeTuaMbBEXZNYAD5KWVcz7rvr3b2Ypqr2eQlbA6tQmikz01A7oag
D8NgrQ9C9OUQbfj9IzM7CYyAPu8R2RAnnzuz2XOotJKIq8P+aslae24uHOrezK5g/WUdzIWhDmJ3
qr7s+WGEnj/mSkT5N8ivEV8kizTviwrc82vQbRmiQ/q466XAaGaoPMoKYOCd50xNuZvhQ4B8yB33
Y1SWSXF2F7A+JP+Ckw+jZsPVCoSh1U7kmhrhTX3iBVXiLXtevW5q/Bl7XZ6VmVvYHoHTeaX8olud
UrObVM7Vv7jYXIYstIj85RsYs3Vslfc4q6P/GBCROe0BjOS2anWpqibntouUFciXnK5U+wXu6ItR
fBn67cxY5Y7qb+JIeSwzvj5MFl/CnZe0Yz5mA0VlvwdM+181ZwrK/zcTV+7AmeqZ/i9P6JFGmdCC
y/JG94UJ7Fxb+JcbZY07lcijlaCUghDc1z2+GMiCbFta9jI9PbBtewYFp8IIIIl08G6lamO3/KB9
CTOeBqFNmsG0xqp/Pa07yqZaLjtByLPet+f5HwXvQS4VgIOIwd+hKDV0Y8OpHbEHqmxEgjpJ8Fmf
epcA1RSFGNTyCcr/YuI2/qlV1ReSg6tSwsBxzdzlj3s08a1hPn7f2eVnAnjL4UVU/llK8IBBmKgJ
p+5btcdmihGWnYqhIoB2nTgoGUVjSjg42rQyvT5/0UrBs9P8d+iIXdSgHDD7yjmrej6ZV6RHzysF
+ybtJgzE+pY0OC8Puxuf2co+I1d8n38fW3/IDAFRoCWxLrw3Ou9TKnqQBEF1s8hwy9LgpF8wW+jj
Vbifrz+OmA8TQJBQt6aiVJ5mjvn7oYq+h+u0NqZAoxNqc7y95CJ3xdYT3cRWJfQFeVBhLqth1IK2
2uBL3rElhjIZDuomfzmXKQbPFScFoXIh1ROpJlupcxYbM57CSzGsYN61zlJFg3aoV21dq04JvH6V
raOgmMNhxcZ3Mg4SQj+gqhCcRw2+85L/Ba3k1M8wy1M+mloUAOwZUtyKY3zV4xy/hewTpJ7bZxiS
+60KatptqzP8Dw9BBtTLQPOxssY96qLwNCUZ2E/8lFQV38/9P0RqTjAh57RAE0WD1vA8HPQOgyq4
mFOekhgFT5R/x49EaZGyRtZpJSviKPEYi/eze1TcGlzMndXkgLTw2vdNSWfLGJb1+16fujUcsJMD
RMul/eEwhyRqJVPTB6AylNtH5toNOS2FxncgwXLWRlarUKYQHzee+kuXnmYVXu5jJ8ycrcLeCSB3
pRRaa5TmzjTDRutoEK3J4+RdZax4PTnmw9WDyVdHPq/19sOb/FMFGzOxxeuN95uB4R9vgt+n1jE6
01PibDt6IntrHBQFyQfPaD4n+AxUqGg/HI29TaTIfqmorxNXhtaYfwavpzZZhfhOdDzgfMry5XKW
2QVw6V87/pVJ41j9Rat1VlUkh4ILl1hyfOFyKCrPd8F6TDfuI5b9dNkCUc+bxCwjIWODUlelQrLE
yT/9BsliYRG8oB1eTYiDqkjhPMFuZdLukY9A4SbY/B/xOryujLg7Nygi9Lb8GWjv+lSSr/lnpKvh
zFS7IaOr3a1dF8qwR8iZOLDgRbAJMZ47Klg2QjuioBeNtZtYIRYnndoth+xsK1fn3rwqVN6oRNz5
YVKFrC6dEgH7dvDN1rDmj/PGNcyOcMElKA+BqReP5wMo9RO7jb0N+D7LQ9eZFY1W/5p3Y67DtMfl
jT6kXJYGbTuzv30A8dd31VgDpEqnnUX8rcrW6oICMcstt3jaL4k4VBqwCF0VWVxu423rXFf72ACd
hSHQbh+6DAqWIp7qtoT5NfJ4OMG9zAJym0ovxqCRmRdeAQ3aEK+PXWlnwrWxshb6ScQ5f6cQQQ91
aqG87khWRzx2115alRBPo21xnnAbAkvA57UjqWwn9UXLvHDECEcryifCirtaSVerlCes/bkKvPEy
yK406WWOz7Xv6ALv1/7HJe62lZbj5QyWQz4TzOWHMWUthbTllYSVycROkLJ3Lz2pid8sivZC4HTm
y4F8LaXKNfXO19tcuVbOQE0/2dzMLbfm7qCMNWrNODgAw/TaE2ldlYED8xaQaGemKfLmgDkd7Q57
xn4+KzMb+TVZ/k8SCnK12UuzQWJGbV/2fAKAdOaLldKAOlFlsb8DZkty8VeBmW8Brupp+Gae5BnH
6j7HkVjWWIIIQaWQhlLXraEMxh/IFrzeGNsG7A4k6uJkT7q3zC9EGIjMvid4JUEQ8QWyLZMoWk+m
yZNdLR26miKD+c/j+GA+snsTSN9jk2rUUvci/6bnMZIsHz7QCdKJMkiSWpWAFJlP8zJ18fRzqtln
YB+a8xUHJ9NPjRlYMCYnRhEVI8iqCdM5tHBSTOFsBJT/Ah3QFm4IAE8a4ACROn45MyHhvy028Uqz
AoKDBAnED9pyGSW4PtuM92v4/7qdvoM57Izn3fGsptR9n0D1UWOlmW1sCSvw9oTvvduLa8njT9IV
sGoIBuOHkkyGxVyVuaSEeqdZ2jw/FQD6zf9ezh9INu+U2PwjTLYGI0JSs5RuNPiDD1JRm6Zw8xfY
blPGjQGFE6mmev9IzUWlKwi4zjA5SrfSQKXqnScyO/SB4dW6UM/Br9X4DEzDSEtollE8U5tE472J
murAnk79PLu4Xcia5bQZPutdLUMXn0lMZ3rCM2ynDMhjec8HKYL30zTBBPkjDEhbnAu8zknOH9GY
qacvWJYXTjFKSTZV9BZYKIYgr8ZFfqK9bx8cCpA51WmZeX88zZiX5Zk6b/eO9452pLVS/2wp3ucb
vN3U01aykKJFZ+ab9qY3nwz7FP+7LVOVy0xJm3jzcBFHzBU6ggOooF476duEoB1uLFOpHgDKIkR2
Ul3OucR5dMkvtUz2les13Oy3vTnQiGa6uMt1COz1HLlb6QtU7xFORVAVcMJglmc/xwj655dbxETy
kjxPtzWyIhqAmcFJxEIk8DiUQVnZc14HxHjh286R8AaLuDKbE+R/LsMMmoVRb/Ir61nN7aazPzPL
D1riTB2k+3h5LAHwIqUy5dl1Eavgp8ZWqBrjAyUYi/5+m7JRIu6sLekDbu5M7V0M0OqjTl9D3Cul
vxzpyhg2S2mJK2Zg3XND2ZOylDug91XxMTDTVZ3FSypPPbSjlL3/Cuhl1FJDXhsslCiiwMXQdahj
43dfg8X1ycDkU5TG3BGf+EDknmMg411apVCTeL4uvb1LhHJzaOhDmLQA5J2NVY890y1xstsb0STx
i5HTFw80YvRITUI3/HWbMqtsyELrsPebxXDILbTxgr4F0o7KN/qjumOFNZSnEK3n1UFCzlIsdION
1MkqYDjJmFa2er1aBXiDtQKTEBSSsbufaB4DipXV+B5Wf+kA6AmlmIiRzsPH5sxeUmjazqcuQrJy
A2GQTdi5/8KoTGziEY1+/PtTMTk30rGUMhXwhh/IcEb6DmPudzdCHDbnYUYSKCl5idOq/YCzkN6p
s0D5tl6CSYl6gv7/U7v0ALo1UXiETAW5Q4wSevQ39yCm4jGjrAo60RE7Eqmh/Q050shzCUtGS84q
mJlTMIZu3nK5WNf+M889mNaEExL6q7JXS58iuLrYZcGGb+ePr0wuHkchxQfH68SbP95Naw50fjih
GHYyiZbc1CYJW/ISEQeyTy7u/ZvNZVXLCzv7b5zegHuh2fccz9THX+tg9R/d+VDR1c5RAZuKBQG7
QmovpFDNTtL2Oaas4KV6j7DMQHqFJXNxkPgY5N+parasQI73k0ne/L6LWEoIHyQk6S7+cbPxPZ/I
20WzV2eKK6ZWAiZKFhBThC3qemM7KeyelksWkrgukcxZXcmhRaIrzM0wfUi0bOctYyJp8mKjQRpA
6dztfZufLRkKaWCupODgxZUYVKJRskyro+FcCMe0vX1EzG0BuL6YiGTxm2U+smrU1f7fBwYVKYDq
shVTj5LlL8stN8t8IGWZSl3ke8fEKnBsREzVMoLkwEnpLa8L8KjSp3gBpbRXHVH7SDSIzTJPWrMq
KjVmXE+LKAOhsquAGSrCkemCSYWaaoNc/FtwHIFyi9/9ktdIwNy5BFVYcIZ0XDxJ224hKgeofa3Y
0c5KeOl+PekZAWgdAzvI28QwdVKrLf3UzcT9v1sRwzK9otrBoUr+Pe5uLygOJ0xBu3E3MYaCWAMd
x31RnNigSuTOjPrsKFgbtfl5vJY/X5hcKduTdlgmya9/ObHFIu2oJU9WpSJdEOjzMDqQBgMihNSI
vUdvt9MNAqqVogfEIkenowXGFuQm63nC3mL4FHgZKuRori2oynl+jQGCv4X79gmgBMal1CUWljXX
U3O7AOS45PBAopzRmMnjiBzbzUM6hYUBn8RLbxmAEeq3plw6aN3E4t/INQcFfYaUotuBvrGtTTE3
EG/qELQIYFSeltaijB3//Qg8PlicuBk9GqxXy9IWOn1T36vHNaJLQMM0SqbrEXZFzyXK6tKUvAK/
V8HSosn6RFLdHJyYquNwpAuRWXhkwYc+1NpruwYNcXlviamZ1qbSmQWLnG/LSoNpavukdc/R8rBv
RxZ6Pb/sGQRdhF2iiBK3kAUv06UEqr0arMRx08VqUbXLZF2Ahbk+317SHvb4a4AWcpmLxVdAxBUK
HiG0OX68/0WgsOXmsGnGXyPrbDGM0cxzAvMgK6FlRgwcgBygVNurqJAM/E5jjNCERRQGa757naLx
T2Y0y6gLau4GjeL5ecYl9GpZW+9aeYizpEjLqr/qlNcqC22oub8E2u/UwvBswVZ52VgBG648JPrb
tbaeyVKCFMuQ+FwQ8T7DP/gLNaq+rGQQhl/rA5akZE2A+ZIh8XppbKhMlWM9Za5MVrHPsP9oxvWx
XiucOINJSD9lazpTXEeJ+tnCiUvzZmRM4CSXR+jErYSzK1xCkOFz0Dvx64RQHILnJGSrOf7KEiQ3
qMUDG+1EkDoCw5mkFFC+liT+j6CHMPxMEz+pKsjs4QmTqqYuVkkLkzmISvDJ6jXdg7I0S/FB60j/
Icn/SmdNsGvsitG8v8JO9e6MwmIl7baqlp3PxhcGG+YDKsjbwOTSh+5vgv5HFPj5VhMa7nPQgs7Y
O3Qn5CcMnLhTH/1yNdibaTwzXUo67Z8kV7LVK80voJEphld8lFfapIJ+wgFrX8crVLu+NRNHvjad
tcX+dMLejJRF8W/NnsCupeiIqDnIpRJf19jMhRLus20hM/dBZ8J19i+MBtY7+8QmhRCwAAqYnG9T
05wm6wFuBzEpirND3A+UhxyYx9sbrW011FC8Y2dSk3vzY/OmuRZ67TzjDXLZsMIA1qUY4wX6ZidE
CPvxkq8C4vvDax0/nIW1pe2x4B/f5Y7ejv+Pj61kR9mTGCdrUtbY71715pNOpspt0wQbT/cB25DQ
vdwtqwHncjEMp2I+vo7Rm5Aw/24GAVYW8FBjAFTR479ocCIj8MKNZpeKiAsT9OCK9ceEIYo20Dff
QEEtGgMoJ1ILcDUcZxCJUowhkzHr7Wo3dQiJOBltHmEteZ7oGD94JQZzkmO/3KUl+L/dj1GLwZxb
UCX2cs04ELYSFdNV2nL/GtzT8eTFhjKtoTma31dkvt5HIkCIL05EAvIYjiGw2AcocpDphwpQBu8G
eaL0jSDdSAW3POYYfNPlyYxsOnwiODsueWLDVasnwZpGxNLFkudLfS9N3ylLxFtgZzTy5Sxx569L
O+ZbEq4wIqQ3oRGoL5Ex0rCX1uK8U0nZsktufa5ly7lQYqA6tyxMLZPmNQt8TvGQOtKPOWm2qpsK
T4qzkTrQeGXEYPg6AOTNDygVjoz9gugzWY5/MwkqhC+Wr4JgIdbhbiEUHgijefjoj5Bxqf15DwMD
qUimQ0QQ8Pz+KC2xW8eFEZfSyxbK0VBPcieChNMit0zRZfK/U1XRy0HsgWW45WwktrMbJKTzQOv/
5ffHIMJOV5ig3CopHSHVMYKVaUZpSocxDU4c2PXrPbx9zrC8oSw3HGvQzRFPDG2xkPcVjynvx0b7
N4gycvZTQTJHhV9yAwgHbIEBOm3rYsM2kd1o6LvibuOYBwlduVhHnt/DDSXV/RN3hBKaVn3EODz2
SEO1Awknt2dz/k6T9cZWzZRT8waSn3BmwYLczY1nTAj42d7tGNVGMyRir/3ReKl12Vpwt47TwOHS
nT519iCs6t7MvXwTzaXkSizJHbrFlQdrqk2ndpGFoE/sVUrYHQG3h/DjTxfrSg1q/+VvadXhbMC7
YYT0ZMGlx7rLO7qOFeeGMviiQ5wi5o0oIFvlejF3WftiU41TRpfrQOKxNSfA881bT8Xgl3Qa9YBJ
eTyIzoTIfsaFoFo75/n5hl3eyz4xijuZ7ywFPX7JvE3/1rWifd9E2mNu3ibtnOtb6Et0kZI8UVdE
5AngymSM3oksOLR0FYnbSHuI72Y2AbyXb9MMxoxeXf+wAZbz/9kshECc+aK2BRFawdSdDEMjnzLF
3D6R14JrtMW6C/vPq+XPvyHHFCfKpx1eyW3CsVOu6KC9fp+duoKNaeKd3sUyYEwQ0bCyMIeQGAB6
6F3xEza+2by4tIkB/SbKKSrxTqhxplZQEN/5nnYzManPIySdJumAaN+vmjummYev4SpPzU0XIglK
xvIUYnpP6ZbHB05X7MBuce44D252dWbfOtAlT6BUCMOXg89CIbbfNpZYOHYr+gMaVWLox/d7H2YG
mu+ic+JKu8tkFFXiMqaxHqu6dKQD6Y8UgbNeAXiPtrNlYVcE9iAQIAIZI3Tg1g3Q7KZD8FryKiLT
GowwKrNtp8Mei0zRLtC0+VOU6PKwWCtYpbs7N/ZWWndJ1IOmM0DFE7tDdahOw6yQgdlJCIb+5yA6
n8TYHtMlM3zQ4ycUvOL+cqn8q0+0kKG5DV/OLuUlVITacc9f8itVRggfAFW0xBRe1y6zrQttOO+S
gzbJ1PQoZJ0Ak1RrT8AVBfmbDuIQa/UdlZdhnJg0+Z+JFxALhA1pJbYg9gA5hnKbNCNJz4+UNxrP
39RXcnCStQ9zz7x1dzKhkzRDBgMBxC1grQVxcDHvGOtPjKF1+2i5+ZT9GESuMMwzYvaeaF7oGLww
7bfsFGBzpjSFUOrGG7CuH0Vu6qQb4RVYmRGzjQTXQEvUJ/yN8TmWgRzSh4o+x34qCvQ8oLwqILZY
EFE/2iZ3BE8yQP0YVwPOPxRIpIVa+r6E+tqw568EPeyZGYl99ItElHsTL9rYiLpMMBxZDggEAiPQ
CYbaZ5YbAhS8tolhLe3W3UR8gLSrOFsATwe+XZUg3bSRwn14PIe3r3LIEWdz1OqHmgU2cdO09eO2
6LvRafLcvHl+J37xhjYJsPcALyU1V94mi7IYr/XelrJD15kzq1onM6oRLjeHpdwtig0X3Mdnh4Zi
ONVxaSd8gX0CZbXJ0WBYuJS2IUsusHB1MJ2yQdbyd69df1Ie9+Y/tkfJ4Y68t6vntjAaBaGgz/pI
SjOLmbJepE75ziB90V8Z8n7y1NhZSBAQ/TKBY98eoBHViQBLkFFFU9yjmMla/mpJB4S7Ojdt6SmI
f2A1VMLwPp78HXpdexKSrdJtaNAVHRW4ExOsbX/CAy0hO+/dX8NHVj/5bZ7HiTbNPJ4z7EMdVi1T
75fv+ZryP9lhuvpgSjaXUpRnu8vb7A/bobcNAr60ACwdrFZSkk26SkZMKTC6/lmy6w1x7Z64Qdxn
Jor0ECpIbMDcjbpRAhgkmJn1pvzrfPSirXMuTCSmciJO0/XYlSXymSRrQkWDx9FR0kMBlsfLD/35
KPbsKl8tji+XZyUWX45XoGdbQQnUczahKHTYWpN1SYutP8UBJJZSx1+T4OeyBjq/KNKUE6Ia4jUX
ACUiIYegv5UBfA3dP63Bfl9+WxF0HGqqtMqWp7nFLgtR9xnfOWivm3DFcgkASqs1N+NH32FpusUO
QGw0HfbSYyOh5CSPM5uzdLehH2PyG9O3t2SJfXXwtzo6BgvcRe7ExZ6xlYOt0v84MH3Sztu0OSQl
SGz65AqGsFIrHw2DcJHHbwj4eSLzSsmjdDxgOzW/efXtp4R2pbib721jl1PvwNejG1ZBvY5ESItH
qpCn9d8CLEBXvSbDsbgT+9NPkpvY8IzJpuWoTY3V9to0MFuHF3D+HfNXo3hI+CNfq+DfK2vZq5J4
Wresa/qp+fhbIe13lQvAwh5dIFljchyMcySUbMqo1pJWVd+u/kzF+94R1O+h34UeOmPyPNoqDxmd
Fk3cX0gilvC5JtFilYnKAmPaJYvs7Mwj9S/OfacTwT8mcsyx31Lh4cgH2PnO3UPgg7pyDCe/JSsx
gWW6T5Nwo8hSG3EaG3HzEVnJ8p8ePrPKpfnBFweBXNGs3wptObtUbkNGjipf8BugeqeKK/HoQk3p
D/MD/81BJEjYDzs8NdEGa6PRwMGYQfc1VLxbB5yWN5qeZ2Mf8VPSDPLA+RdV/ADmM0r1TTtKO9GM
zCVgfQqe9Qc+1eAsKMq64jovV4iH2GcMAi+wyx3RzFVAwrMI6//0qqr+ukqQJmcmJ8ZsRekKiDor
x9Jw+H1niGOvEkAZef6R0bvkJeiG9oNqSuY+v+q+9gUlGvr2HmUZqwvjFtv1133WQbbA4C8kNodW
ELgkzWbnMQx4Yc1x6DgM3kHstfbwPqfZXbjn1dFXSgLzQhB8ABGrY5089PHXwP03SV8bUSOdskzL
3QIjmkmAj/cy46WhQE8Lny9qWWB5cL9cBJ2stpOXseXpl+2pochCz9J5i9jdQNQ2oxGtqn3YddLH
9190Swt/AZI66hlQwHGFJJULqS2VGjgbTlS8OccYpTNQYbAg808+GV+YoRKOMcKUcbyCY8gM5hmD
86PoTYZJsWBd152C5r6yiJ1Ma6G8KYsGtV38yPhCheOrbwDK2fOEC8zpJOHvMZ0tfxPgYmr54cQS
c8sUAqhjPwLdUka1C6GZmjNQhfTtL6ctensq2tPQ8VFe/yy0rbRH9aTPog4pnNb/dpNDbYl7KN0q
XiDXl2xYiK13LZT0et48263VEnBzGPZlyfPLHIc4DrOx78jSz1uBykhKUC9y14iIiTi0vTdhHjhm
WGMtX4pHwYd5/lYI1kCDZFwp51tb7eTBkoUSJuVgubgMqT1b2gNKLp18f7ulu5MlP0VW1JRR4Wef
otFCLECoGF6IfGGizuc7mlxEBXmbfOW4JGydex4J4Q2l1jLDOOY0X5Z7zk/e8b4U/vyyDisBX1ts
NVckNd+l5dQABfWn4jt6x9DzW+RfmnUf5f41ZXLJ1koXYojrxuDXd9lCW4La9m3M8n9NVkn05XOU
oKGxPwM4fiwYzdXCbLVxEZHeC8najZa6xkmIqipy8R5/ZoURv0gsRPtTZsayZDN+d4v2gUm0qh6i
zn34aMrUGf8UClYgxvqEONOiFN42qE7GFArykeB/GOfafRUivitWAJRaKcF66EsFjjliz3gBq5vX
dpRPZTHyYHMbl7T5+VDQYQzVtgoxvoZ3oa3BDjiN/ehcizAnp/qWENPWIpw0z8f0j63bvXgO7JdW
bginetCiNRB5tMBqFX/8i4gG3MVf/6xW0itJtBLFUNqGUTOJdaZuMZwSUpsWAzIiXvf6BQn3FNTB
1xZgJ5LyiIDYtflkw6qwyLaZ25rGC97BSUbViHCSNsAao4y2abD2sbeZMSC3QLrpwHnTkd37EsfQ
D46zN6KHWPZ/1Up3nZHvVDm3siQvZnsTlLLkq1iXP5xQ8+n02GTO0F2WshOZ2Tl38avGN5nGMEwj
EGGZbce8H/gT8Dk3YJhbDp//nR5JFGcRAjxUzM1X0liThgJckWyIoB1i12aaGoQB+Qb4Q+lzVaKl
9Sp4L8xFOxKFA/aeKWY3hnMpxHgXH2gacuddDY73P79+HzeRO+1Tk57gDjL4n37LGLaLvVi86S2Q
LKhyHRZYN76+amQbvNNuXCN7F0YifBgqEeB3Ih9KVjpm9bYXX/El68BsIXtHgPLoiB/HvRSm9vk0
OZhUG6q/5xI6q/NrOB2gjZm4p/4Clne//16/hLijU1SZCno0B072CcayLDGg9t2CGJVq5g/S0YTR
eck5bfJj4i5FCUN8FgmDIoeoE13c/oZvbJo5FXtI2DiXk4lET62G9VpNlQx1RYncZ9KOB3l9ktAg
v2Lfqwyzh9bxANzT75wAXHPerdHj2kBe3t9nLB0/8tLGF5nVRW4uvXNrTn7JQjuplXgCDLs6vw+2
nyAQ5dDYssADDtWYr1p+6RWlkGLI9PTNAEDah5hrAmi9ApWELUENvRzS3y1CDLwGqrqlMmh8wPSM
blBeZhfF5/DfPF+RVpYw+ddZkqHCWyJc6xlC5X2LkG03FKe45GqmvwffoKzdRVgDYqQNs4v9vKrG
E7DCq0pWeD8djFsAzIF8ba4ScXitCtBcCyXsUy6foqqhH1lbnEEATN65uWACtyku4iK8xbbiZCuZ
rKj8bEobVJ8eZJ5fSqJL04ve0yGi88sUSGcTa2Vt9y1R0XowrkPYWCFAMPAA88f7Bm5O/k/+L3WJ
75Ss4Lg6aSIesq3/DzY8GBlnAeCdRLChEyvfMHW3HpCcrjSTGapMCGgPpCXYFujCN2eM9aDiwaZY
Qi8FeP3qdmrZUn6nlJU0x3pw+u48L3FyjUBcdlwkNDluJan7MpiWeOGXwUkgmdkAeaxINNdkLZzs
bSE/u7J1MjEcEam6kZgb2V7d9sTKuze6ITCEPCpEGpsSHg7KZQuIpEP51UI+v/K7KsOQaVLy41ID
q7eQpu9DJA0PWxb8Mmgu02OAQWTijhFOHBkAdHXLu6Qpy9Vr5rc1XxPGZVaSCPS2Ys77xkSJWCzS
/BP1cdBZ4e8fWm9/iX+mK5H508B931kgAKhjXytUvI2dup0yzdWrk+iIH7arCGsls1t70zb2ssfk
XbjGtMneCQv6AYBpmg3JU2ntN7tx66LMCDaNAIdyft/0XmNxasUaVuySprGdpf+67/kAwg8d+OSz
2moEphnMYG8dpyQe39pJrYbb23cVJxRCrrBK8Y1NyWp/YdYr9FcWtkQRz7F27l+h50kJ0BfT03Q+
UvRi/TkAlok6dcky+5hN8TrZLGMUYP214reEWZaUkruOECfbn2/S4va3sz7N8nbL2NBK/0hxvxQs
gJijmEBudBWjvo5POR/Ge5jTO1WHlMfmvJInYh5qYX3VaJu/0KqyFJcQOIAaiC1Cco+b070zLhn2
yf/vXPYo8neDRI3YJ6ZDV1yfU4twE3IKS9ohxeZB3qBINda5sSXLAxMRpQFiW+SWtNGKP2WoFhWC
HRro3ZVRB//bRCbVxbU0mXFg6MD/RaQGyCz9RCj8cdLbPQZ0ViO0xcJHw5aUBkX5NYHv40iP5Eq6
l/79FuvzZPJXldxqjmrFMCFykN5Z2yYfEc0fTzHBjp3znkDY/si+5PU1YedHczo5tKd3HZ1jv3eA
O/ci4yiqEgkfRUeMWyPuMU9OHKlVka392QvTvwOkuOly9jvAcOnIOZkyC1s6rQPHsSpoidHUp/Eq
l3icGAIsiXnn8mslND5u1DJu3riMp04nF1z3MZqejGcKrtw+qUczOxOxhV4H3vrDJ0coRpU69/45
S0YRE2fwz7IfevlJ47e9yj3q8khk3CWCWAXW9Poea7EBPiAodGujybT+/hsUjxx23MV1YDoEWpGb
OjM6YJ++HpI1pvjz623H797GxDYh1jf6V7yPBK1nPYdNop2IpbWdKPnHLIH7g2iKvd1CCcFT0GTT
TcgCsZcb0cRTJlgh1x47VabEwP8NS18SNLhAMZ2lz2iwTkIQdQFtA6pr9jjwk+2lbBN8sw3xqGYX
nyGuOtQIGTOOU1rTN9/nzyeE/VPMPSe7/yb38TyRLD9UZtT5pKhO7M5Jr30nvPe7bUcZc2UP4i51
6oczdvAf6qWn93XkM7mK0117d0GL4Ex2+1jsabxUPSKlOmiYFkD/58Z2iThs+y3BxyxV6GCQPtQp
+JiSGVodtClHyYRZB/77NS0UV/nQFJUhaq1nqb7VK4c/GezH2ihLMpi2dFc8N5cWW8ad5FIU3u0M
JmaOdQwobN1zkjARn17oOkNT16rqirfXuoSMr16ownnEqLs0glsGE4WOFToDDSWxCMtDj5E5u4o4
03mkxvZU8xbGzpPQaccn0vNERHIoporzNpY/TZtwlFEdzjtN9bHkxh56cYIbh7Op7gWCy5VJfq+X
8UDXG8SALJ7/v+RBfbmTdYbiG6nJjCpswbIvHrUuPBnlFaXB8mvgfYVKNAlka1bufRJU1cFaeVi0
ZKJVlRsySbfbGdNRQ7N4kb9EfoIFUXmPVydkL7SnqSi2oyRI5Fn+gYR79QCTMHuaFYAss47dUvRa
bcp7BcIv6k3rh7BC7MG77CAQJwybw3F52kvLe2fHnR3fQ6Kt8mWMy7Za1WvxyDeH7W09t3qlWYL+
65AKQg0lLavvVpggEIn5YmGHZOT+wGscUffWjhaxyVUsB2iSL01TfFerYpYEheKg3z9KQZ7Fj6zE
ukLls3mUJjqL7jxu6BD347t4NJ8sTbl7Fdjz8K1KQbYBILCSyeBD+ga5iOXGlzxu2zs9aOzB/iix
RRnqeGU/OxpijnyqkiPVJlIEaiEp+Z8JNmcZzPJqf5ockU2SfVCK+KsNBqIkt0zuiAPfcaPEzagA
goJCgqTR3RlSfdgt0/SG4A3sQ54GYvXWaD57XsNlW1Xb//BYlGy6Q0V3RiGa+qzxVNCSVprsCZqT
+5Ac58AiFb+z195Zht/9pe4dOouhDi0LvjrAZr3RuzHuwpC+kE9h7d+V65kZYevQfyOSqQ+sJTHR
GRXGcBfmu51K+JIWgjtuBuY0LzBJ+EErwGwj/2AldRb4Bh9PlZczZLLWT+HhvMJubPd7vY64Pzmg
5Js+b1/afkSsbVMbrkPONuDkfkBeLTtRpcNn7CMwGmXAngA7GXPdfzXK6JxLgBW9/DGp3NrmFW2Y
/raUk/vcG0Tja0FthiacBahjB+LziPuFv7iiMnZAtma+S9/MFeF0w8CYQZWYL/e80rFH0Lt9vDlc
R7DkxwmHk9vkmF9hSOeg3RAt7aP9D5vxok771YLnczjpFwbh4TAUUkxXHMmx77MCxk71B1vzVny3
b4mkqTGtD4KVyFae/3MpZ9gOy7r1nWoBzbcUI3QTZ9LxQsiNUxNQWjtKx5O8B7b8pxqia8teP2qL
9SOX8PIxCZWvxOvUhUF7wga2LF/htFwTBjxpAfdt3+jkPCsKnmak33ZjVR26G16dTEfct8B+F2Pn
VnZR3yJ/T3+WnrhO5QHFVVzN6EOlJgpgBy0xFiDPaRwZoSo3yWPhzLPOZkyDhtwo9pXqxWOzNtoP
hCforEp7EwYIHFHsFFb4KbeolZe7RdRiTPP3Z56lx3ynq70PbJhkSYUlRnlTV9p95a3bp8RhDhPR
+8swd9SsHG9MyXlHJWIXW53CcjsOIxtVbhnRDNba2QSKKbwPX07ygPFITk28cV7RIrOUAYwH3fri
jhvG8sioFi2QIAXBtDnrGoGk/KJSFwRp3a0ai7JOQmmgHYgVQZNaYOeD8r3uHoKVI38eWGhh7Bja
3sBMPITO+UJ3E9e0N4yWBp4qSnjVq8yNQxddBS0NDJS9y7BMk03fneiXsNvmd/23mzV2YfiiYGhL
u9lVBU+06bdQr9CQ7WBvQfM2nxuKsyTgzWzBB1xOKUrGIa4vPbiScVIYxpfOK/2gKOEtr/FnE8gj
NO/KGv1OUZPdcLbRJgw8u0f+Wb1v5AUJWX9KLXDntRuN+GhxwRPD5wmcM3pMx9HuwWo1EThH3We9
SQiy3EaiS5EwU+pzhlIpN2Qtc+jpeEhtOQ6CoZRKa/ILHLf0jaknhhAyB5QJvGvmOyGhE3fibFwu
aThgjCet3DZ3RybmkWFo8iVluo84hnD491HK0UFSGblahbiPqXgkJeK6ZUp5oNa8zOKceTLmjhT6
3Iad78ke9MwdF21liYBfGFDpqv9MpAlJld1UKt7UnF22Gzlqzwy09cbILMTwHTrf9Ij8BrYFoAZw
GMO4QQFMhiqT4v3N9XTuEv19oF0ZE5D+Zf1YkvR8rQqEM0XiPrZphokVFG3dmgr6M9G2vmXnf3Yr
hrA36BfrlPeqdmX9vrLKDQOtp1v17rHC6DkAgwXExS7fbjh1UHPFeP+NPvA/4tlacVGreCwcxpm+
pibOSPxL4GD0XujaghF356vcrNHdR4ZZddyKz6fA8cCZ+ducbQo1lsA0jtQDW9fWIQf4jrRC6adf
+LW6RmMlG10n/su4MmxWb/ujeRiXzr0cuSxywFYuiiddxJpVXnrQnvC6nkHmevHc+xPyWcxSpgP5
mnP8ktOxZwCus4TH0n8PGeUYNig/2/Vp8ssvYDxuWT4qmv5EHnMJrnry2BcKY2Ibkmm6H+KWJTH6
OwtpVR7LRwQ3sDjXEspp9PgdPPTGOSxvoSms61PUd/OX4sIuttHG2pCaITIxmr6n4Nth3F+Rg4mk
P04uulizL0yzrJ7kgTjr3s3XSStHFC6E/bYnke+4yOuQGfqFqm7Sm4vNEfUbvSrCN70M1d9BWB46
wfSIPEWu28GKMJJO5DwoDQ1k55vqlGYs1eIiWqHyNEu2pMy0rvtF2jP1E+TO7HsuxYOQtFp51Tcj
IAugWraJcXQsocdKrk/i9Noe5vXLxPfoBd8kr+T+0NLTw4mlJXv7Xps+fm6N0NWeOgBAJDT8V9KY
0sm2PkXquJHDvXcCrAlydtHnjuVpqCcG6Fw5xNMnDBXCcpgEG85a/4NIr2oyb0r2JmkY8MOJpkrU
INFs6MDR+sh1lWzzswZTof5vznoAPxj3rCiOXs4QbMoSdX97mYc7z6DpuYAR/zy7j1ZjqpjyIJBV
LyT8F9ZSEvFOgL5Bs53sDX/bGvDQpTgz8nFrd5FtXs5yXgoc8EQyZXjCeR8ONOgpBFrzWJw+vy0J
V8Os1NxuWp3laO1GA/P/j/AClFeqY8QCpnpMtzEMushRdkkAkZARe9wwsFQjlv/6/hrsfE2KzGee
0zqrRnXCRIIuTheT8YTk86sr4sqp+yHpEZzRcSKjs8wRGvUEG8sdmsGJUDjz9g/UhJye/tZ5lD3+
UK5E/Y5wqKUrN0Lsu5A4bsU2YBALJSXuXiS9I89v/RB17HpvVq0noDoAHJtIMOFdFX4CbJ7RMUHc
dcWYR+ixSBI2R074jw6ZKSdnulniWxAZxqGPQCV7/zeajpTH7xVcFMGLQ8TcskzxWDeNgVQm3z9h
GEbWZxgtaOtZmmEQZE5ar2I2ZFsUUAIFq/NabyzmF+6UbqcwaIP/XeNa3Xct96+vBxkEzuYxFxKD
YEqvWxmF9/XHGf1iUwWB9JONNQm60XCxL+j2rd45PghpvbDCS2jCxzJnYYcSoC6UH1hsW1UidlrI
33wsf6AXyWdwAqI0B200wEyP8IUb5q9cllgRncMAGF4d6LP0BwD24Ao/QH/I2BjNjTGQzHNmDg0N
kdDP5lyVmURJY1l1IvslP4T9DtKhRUUKmH/sTOeRW9Ta1J0AvrBg80WL0A1roWdQ/4bei+keqQyA
rdDQtI1UYURLjIt7MtvEPcOAzuxWpnCvff/g2eqtJhuOukGdWxfDoYzkVn9uJY2w8QId+ZBnA4eY
OAs+hLFV2zKbL164NOcJpfNQnyamsaJruE9UNCPHynVCa+BUT1uF0qQN8cdJR9lJiySpQj9hwROM
+EU+dBE0r5dJfQ3x3etv5seS03oiKuDy1g4xiSRVWdubHiVbgbmnzf4nfw7K5EQhRxtOa26ubqkY
teD44r3l3pRIPh+OzQ0sF2RWOe/X1jye2GjcNUK3b20JcjM47hw9xpgxoVaBN9yumQCKb6BLvse9
/dyd2Xqf0Gn2vLfHku2n3kEU8bp6ikfayVgYA8DkWemM7Kh8GgGdRj21yJ2ZmzsuVXIQsRpEso++
spGF5uezJn5w3apnKd/fYMm41dte3eRZ/N0Rv0MU6Rztpfp8vb1E3CRWu0hQGBSus9gbYGsMk1S0
syI4N1sPXY+OJ+ATrh0ymJGYlURoPhE+wYCHkAOpyt4zN+AtjPc0jKTymOxfsF8+rhja5VxDhyY4
5E8cqaJp1RDfpJs+9N0uR1wm5EfSFjLJveI4sXvF9XPdOotyAp5Q8bJ/gLQ3TXpwb8pJSqXNQ76+
KptBuJCjSM8S8VntY13cai5MMu55rO4HqEfxRp8jQ1Eo8hDYsQ5GtHqIflzOy+K5juPT5kC4XbVK
HwcS07Ij0kxmNGxpxZLe9tuOaAPpGVEEmc48SJ4ch8wNudIlMNe45SgrBPvKsqw7jcM0W638OhCS
fok8pd4el1GeTfhASgiTWk8r2wsfi9fFCjgY6p/gtYWXQLrsXe2xVu6V4NkCEtzvwchpwc/MZYRR
OiioxyE+vuvTSvY1BVFzWd/EsQDb6jmE0kiUw1eJiAvtM172aDN1sJoNa4Tne4/G2FlmEUwtmvmp
kW+FD0U9hyEzbXSJMCyN5113STxZGRoatAsUbt8wdEBw+1nbYOjQy9YUtjcnd6HAYRCTOoYlaJZo
jbLZTW57LG2EYwRyGxgTdKEgIvmjWUH0/L8kZhgerq/ILalnBppwWiOgz4OARG8vYU1pJPMYnfZs
3y1KQcWXY4D6CROQcYdtq8mOYt4bMfIFXQp4FlhBzlqtz2Y4aiQny2qNYSWX/M6XSK+Y9pyTIlqr
3llqUD15UrgYIbA0zHbi5h2WIC3oxfmsProzkvT0s7VYbHQvnyO0TRvBNZE3xMST5vWW+9y0KPyF
e/dkjXmvosuq//jaynv7do86RgEfsfOhSKzPu4+GnbglVLUJf6Xtrox+h5WDuB+D7TF+urRdxnt9
ifRv3Pnh+XF5Bq4=
`pragma protect end_protected
